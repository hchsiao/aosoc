// Copyright 2017 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the “License”); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

module sp_ram
  #(
    parameter ADDR_WIDTH = 8,
    parameter NUM_WORDS  = 256
  )(
    // Clock and Reset
    input  logic                    clk,

    input  logic                    en_i,
    input  logic [ADDR_WIDTH-1:0]   addr_i,
    input  logic [31:0]             wdata_i,
    output logic [31:0]             rdata_o,
    input  logic                    we_i,
    input  logic [3:0]              be_i
  );

  localparam words = NUM_WORDS/4;

  logic [3:0][7:0] mem[words];
  logic [3:0][7:0] wdata;



  integer i;

  always @(posedge clk)
  begin
    if (en_i && we_i)
    begin
      for (i = 0; i < 4; i++) begin
        if (be_i[i])
          mem[addr_i][i] <= wdata[i];
      end
    end
    // always read data
    rdata_o <= mem[addr_i];
  end
  // seperate to 1 byte writing
  genvar w;
  generate for(w = 0; w < 4; w++)
    begin
      assign wdata[w] = wdata_i[(w+1)*8-1:w*8];
    end
  endgenerate

endmodule
