module M_0
(
  output reg [8-1:0] Q,
  input wire [13-1:0] A,
  input wire cen,
  input wire clk,
  input wire reset

);

  always@(posedge clk) begin
    if(reset) begin
      Q <= 0;
    end
    else if(cen) begin
      case(A)
        //32'd0: Q <= 1;
        13'd0: Q <= 8'h54;
13'd1: Q <= 8'h55;
13'd2: Q <= 8'h00;
13'd3: Q <= 8'h04;
13'd4: Q <= 8'h40;
13'd5: Q <= 8'h54;
13'd6: Q <= 8'h00;
13'd7: Q <= 8'h00;
13'd8: Q <= 8'h4c;
13'd9: Q <= 8'hdd;
13'd10: Q <= 8'h00;
13'd11: Q <= 8'h55;
13'd12: Q <= 8'hd4;
13'd13: Q <= 8'hdd;
13'd14: Q <= 8'h00;
13'd15: Q <= 8'h4c;
13'd16: Q <= 8'h50;
13'd17: Q <= 8'h54;
13'd18: Q <= 8'h00;
13'd19: Q <= 8'h00;
13'd20: Q <= 8'h00;
13'd21: Q <= 8'h40;
13'd22: Q <= 8'h00;
13'd23: Q <= 8'h00;
13'd24: Q <= 8'h54;
13'd25: Q <= 8'hdd;
13'd26: Q <= 8'h00;
13'd27: Q <= 8'hdd;
13'd28: Q <= 8'hc4;
13'd29: Q <= 8'h5d;
13'd30: Q <= 8'h00;
13'd31: Q <= 8'h00;
13'd32: Q <= 8'hbd;
13'd33: Q <= 8'h01;
13'd34: Q <= 8'hbf;
13'd35: Q <= 8'h09;
13'd36: Q <= 8'h9d;
13'd37: Q <= 8'h11;
13'd38: Q <= 8'hdf;
13'd39: Q <= 8'h2d;
13'd40: Q <= 8'h00;
13'd41: Q <= 8'h00;
13'd42: Q <= 8'h99;
13'd43: Q <= 8'h00;
13'd44: Q <= 8'h00;
13'd45: Q <= 8'h00;
13'd46: Q <= 8'h04;
13'd47: Q <= 8'h00;
13'd48: Q <= 8'hfd;
13'd49: Q <= 8'h00;
13'd50: Q <= 8'haa;
13'd51: Q <= 8'h1e;
13'd52: Q <= 8'h08;
13'd53: Q <= 8'h00;
13'd54: Q <= 8'h8a;
13'd55: Q <= 8'h0b;
13'd56: Q <= 8'h00;
13'd57: Q <= 8'h00;
13'd58: Q <= 8'h08;
13'd59: Q <= 8'h00;
13'd60: Q <= 8'h00;
13'd61: Q <= 8'h00;
13'd62: Q <= 8'h00;
13'd63: Q <= 8'h00;
13'd64: Q <= 8'h15;
13'd65: Q <= 8'h3c;
13'd66: Q <= 8'hb1;
13'd67: Q <= 8'h15;
13'd68: Q <= 8'hd4;
13'd69: Q <= 8'h34;
13'd70: Q <= 8'h3d;
13'd71: Q <= 8'h35;
13'd72: Q <= 8'h69;
13'd73: Q <= 8'h77;
13'd74: Q <= 8'hbf;
13'd75: Q <= 8'h4f;
13'd76: Q <= 8'h75;
13'd77: Q <= 8'h0c;
13'd78: Q <= 8'h29;
13'd79: Q <= 8'h08;
13'd80: Q <= 8'h6f;
13'd81: Q <= 8'h7e;
13'd82: Q <= 8'h1a;
13'd83: Q <= 8'hbf;
13'd84: Q <= 8'hfd;
13'd85: Q <= 8'hff;
13'd86: Q <= 8'hff;
13'd87: Q <= 8'h07;
13'd88: Q <= 8'h00;
13'd89: Q <= 8'h14;
13'd90: Q <= 8'h33;
13'd91: Q <= 8'h2c;
13'd92: Q <= 8'h40;
13'd93: Q <= 8'h44;
13'd94: Q <= 8'h18;
13'd95: Q <= 8'h00;
13'd96: Q <= 8'h00;
13'd97: Q <= 8'h00;
13'd98: Q <= 8'h00;
13'd99: Q <= 8'h80;
13'd100: Q <= 8'h00;
13'd101: Q <= 8'h80;
13'd102: Q <= 8'h00;
13'd103: Q <= 8'h8c;
13'd104: Q <= 8'h00;
13'd105: Q <= 8'h00;
13'd106: Q <= 8'h00;
13'd107: Q <= 8'h20;
13'd108: Q <= 8'h00;
13'd109: Q <= 8'h80;
13'd110: Q <= 8'h00;
13'd111: Q <= 8'h80;
13'd112: Q <= 8'hf5;
13'd113: Q <= 8'hfd;
13'd114: Q <= 8'h00;
13'd115: Q <= 8'hd4;
13'd116: Q <= 8'h00;
13'd117: Q <= 8'he0;
13'd118: Q <= 8'hc0;
13'd119: Q <= 8'hc0;
13'd120: Q <= 8'hf4;
13'd121: Q <= 8'hfd;
13'd122: Q <= 8'h80;
13'd123: Q <= 8'hf1;
13'd124: Q <= 8'h80;
13'd125: Q <= 8'h90;
13'd126: Q <= 8'h00;
13'd127: Q <= 8'h80;
13'd128: Q <= 8'h00;
13'd129: Q <= 8'h00;
13'd130: Q <= 8'h00;
13'd131: Q <= 8'h80;
13'd132: Q <= 8'h70;
13'd133: Q <= 8'h40;
13'd134: Q <= 8'h50;
13'd135: Q <= 8'hf0;
13'd136: Q <= 8'h00;
13'd137: Q <= 8'h00;
13'd138: Q <= 8'h00;
13'd139: Q <= 8'h90;
13'd140: Q <= 8'hd0;
13'd141: Q <= 8'hd4;
13'd142: Q <= 8'hd0;
13'd143: Q <= 8'hf0;
13'd144: Q <= 8'h00;
13'd145: Q <= 8'h00;
13'd146: Q <= 8'h00;
13'd147: Q <= 8'h90;
13'd148: Q <= 8'h00;
13'd149: Q <= 8'h88;
13'd150: Q <= 8'h00;
13'd151: Q <= 8'h08;
13'd152: Q <= 8'h00;
13'd153: Q <= 8'h00;
13'd154: Q <= 8'h00;
13'd155: Q <= 8'h10;
13'd156: Q <= 8'h40;
13'd157: Q <= 8'h00;
13'd158: Q <= 8'h40;
13'd159: Q <= 8'hd0;
13'd160: Q <= 8'h3f;
13'd161: Q <= 8'h0b;
13'd162: Q <= 8'hd9;
13'd163: Q <= 8'h05;
13'd164: Q <= 8'h51;
13'd165: Q <= 8'h03;
13'd166: Q <= 8'hfb;
13'd167: Q <= 8'h9f;
13'd168: Q <= 8'h6f;
13'd169: Q <= 8'h25;
13'd170: Q <= 8'h04;
13'd171: Q <= 8'h11;
13'd172: Q <= 8'h0c;
13'd173: Q <= 8'h21;
13'd174: Q <= 8'haa;
13'd175: Q <= 8'h32;
13'd176: Q <= 8'h63;
13'd177: Q <= 8'h03;
13'd178: Q <= 8'h49;
13'd179: Q <= 8'h0b;
13'd180: Q <= 8'h00;
13'd181: Q <= 8'h00;
13'd182: Q <= 8'ha8;
13'd183: Q <= 8'h63;
13'd184: Q <= 8'h06;
13'd185: Q <= 8'h2d;
13'd186: Q <= 8'h09;
13'd187: Q <= 8'h22;
13'd188: Q <= 8'h00;
13'd189: Q <= 8'h00;
13'd190: Q <= 8'h04;
13'd191: Q <= 8'h00;
13'd192: Q <= 8'h0f;
13'd193: Q <= 8'h0d;
13'd194: Q <= 8'h9b;
13'd195: Q <= 8'h2f;
13'd196: Q <= 8'h02;
13'd197: Q <= 8'h00;
13'd198: Q <= 8'h02;
13'd199: Q <= 8'h00;
13'd200: Q <= 8'hee;
13'd201: Q <= 8'hdb;
13'd202: Q <= 8'haf;
13'd203: Q <= 8'hbe;
13'd204: Q <= 8'h08;
13'd205: Q <= 8'h88;
13'd206: Q <= 8'h22;
13'd207: Q <= 8'h0e;
13'd208: Q <= 8'h20;
13'd209: Q <= 8'h00;
13'd210: Q <= 8'h01;
13'd211: Q <= 8'h00;
13'd212: Q <= 8'h00;
13'd213: Q <= 8'h00;
13'd214: Q <= 8'h00;
13'd215: Q <= 8'h00;
13'd216: Q <= 8'hc0;
13'd217: Q <= 8'h00;
13'd218: Q <= 8'heb;
13'd219: Q <= 8'h0c;
13'd220: Q <= 8'h20;
13'd221: Q <= 8'h00;
13'd222: Q <= 8'h20;
13'd223: Q <= 8'h04;
13'd224: Q <= 8'h50;
13'd225: Q <= 8'h54;
13'd226: Q <= 8'h00;
13'd227: Q <= 8'h00;
13'd228: Q <= 8'h44;
13'd229: Q <= 8'h50;
13'd230: Q <= 8'h00;
13'd231: Q <= 8'h00;
13'd232: Q <= 8'h55;
13'd233: Q <= 8'h5d;
13'd234: Q <= 8'h02;
13'd235: Q <= 8'h06;
13'd236: Q <= 8'h5d;
13'd237: Q <= 8'hdd;
13'd238: Q <= 8'h00;
13'd239: Q <= 8'h2c;
13'd240: Q <= 8'h50;
13'd241: Q <= 8'h50;
13'd242: Q <= 8'h00;
13'd243: Q <= 8'h00;
13'd244: Q <= 8'h00;
13'd245: Q <= 8'h90;
13'd246: Q <= 8'h00;
13'd247: Q <= 8'h00;
13'd248: Q <= 8'h55;
13'd249: Q <= 8'h55;
13'd250: Q <= 8'h00;
13'd251: Q <= 8'h09;
13'd252: Q <= 8'h54;
13'd253: Q <= 8'h51;
13'd254: Q <= 8'h00;
13'd255: Q <= 8'h08;
13'd256: Q <= 8'h10;
13'd257: Q <= 8'h10;
13'd258: Q <= 8'h0c;
13'd259: Q <= 8'h11;
13'd260: Q <= 8'h10;
13'd261: Q <= 8'h00;
13'd262: Q <= 8'h11;
13'd263: Q <= 8'hf5;
13'd264: Q <= 8'h35;
13'd265: Q <= 8'h88;
13'd266: Q <= 8'h08;
13'd267: Q <= 8'h10;
13'd268: Q <= 8'h00;
13'd269: Q <= 8'h00;
13'd270: Q <= 8'h1d;
13'd271: Q <= 8'h19;
13'd272: Q <= 8'h80;
13'd273: Q <= 8'h80;
13'd274: Q <= 8'h00;
13'd275: Q <= 8'h18;
13'd276: Q <= 8'h01;
13'd277: Q <= 8'h00;
13'd278: Q <= 8'h02;
13'd279: Q <= 8'hbf;
13'd280: Q <= 8'h08;
13'd281: Q <= 8'h00;
13'd282: Q <= 8'h18;
13'd283: Q <= 8'h11;
13'd284: Q <= 8'h00;
13'd285: Q <= 8'h00;
13'd286: Q <= 8'h00;
13'd287: Q <= 8'h18;
13'd288: Q <= 8'h03;
13'd289: Q <= 8'h3c;
13'd290: Q <= 8'h00;
13'd291: Q <= 8'h03;
13'd292: Q <= 8'h90;
13'd293: Q <= 8'h80;
13'd294: Q <= 8'h21;
13'd295: Q <= 8'hc6;
13'd296: Q <= 8'h03;
13'd297: Q <= 8'h03;
13'd298: Q <= 8'h02;
13'd299: Q <= 8'h03;
13'd300: Q <= 8'h00;
13'd301: Q <= 8'h20;
13'd302: Q <= 8'h13;
13'd303: Q <= 8'h00;
13'd304: Q <= 8'h0a;
13'd305: Q <= 8'h02;
13'd306: Q <= 8'h00;
13'd307: Q <= 8'h08;
13'd308: Q <= 8'h60;
13'd309: Q <= 8'h80;
13'd310: Q <= 8'h00;
13'd311: Q <= 8'h03;
13'd312: Q <= 8'h17;
13'd313: Q <= 8'h00;
13'd314: Q <= 8'h01;
13'd315: Q <= 8'h02;
13'd316: Q <= 8'h00;
13'd317: Q <= 8'h00;
13'd318: Q <= 8'h48;
13'd319: Q <= 8'h0a;
13'd320: Q <= 8'h10;
13'd321: Q <= 8'h01;
13'd322: Q <= 8'h00;
13'd323: Q <= 8'h00;
13'd324: Q <= 8'h10;
13'd325: Q <= 8'h00;
13'd326: Q <= 8'h10;
13'd327: Q <= 8'h08;
13'd328: Q <= 8'h75;
13'd329: Q <= 8'h55;
13'd330: Q <= 8'h10;
13'd331: Q <= 8'h90;
13'd332: Q <= 8'hd9;
13'd333: Q <= 8'h10;
13'd334: Q <= 8'h78;
13'd335: Q <= 8'h7c;
13'd336: Q <= 8'h02;
13'd337: Q <= 8'h01;
13'd338: Q <= 8'h00;
13'd339: Q <= 8'h08;
13'd340: Q <= 8'h10;
13'd341: Q <= 8'h80;
13'd342: Q <= 8'h08;
13'd343: Q <= 8'h80;
13'd344: Q <= 8'hb1;
13'd345: Q <= 8'h8d;
13'd346: Q <= 8'h20;
13'd347: Q <= 8'h01;
13'd348: Q <= 8'hf0;
13'd349: Q <= 8'h18;
13'd350: Q <= 8'hb8;
13'd351: Q <= 8'hbe;
13'd352: Q <= 8'hf8;
13'd353: Q <= 8'h04;
13'd354: Q <= 8'h00;
13'd355: Q <= 8'h00;
13'd356: Q <= 8'h40;
13'd357: Q <= 8'h00;
13'd358: Q <= 8'h80;
13'd359: Q <= 8'h90;
13'd360: Q <= 8'h51;
13'd361: Q <= 8'h00;
13'd362: Q <= 8'h40;
13'd363: Q <= 8'h01;
13'd364: Q <= 8'h00;
13'd365: Q <= 8'h00;
13'd366: Q <= 8'h08;
13'd367: Q <= 8'h04;
13'd368: Q <= 8'hea;
13'd369: Q <= 8'h80;
13'd370: Q <= 8'h00;
13'd371: Q <= 8'h08;
13'd372: Q <= 8'h88;
13'd373: Q <= 8'h08;
13'd374: Q <= 8'h80;
13'd375: Q <= 8'h88;
13'd376: Q <= 8'hf9;
13'd377: Q <= 8'h00;
13'd378: Q <= 8'h00;
13'd379: Q <= 8'h00;
13'd380: Q <= 8'h00;
13'd381: Q <= 8'h04;
13'd382: Q <= 8'h00;
13'd383: Q <= 8'h09;
13'd384: Q <= 8'haf;
13'd385: Q <= 8'h1a;
13'd386: Q <= 8'hbf;
13'd387: Q <= 8'h33;
13'd388: Q <= 8'h15;
13'd389: Q <= 8'h08;
13'd390: Q <= 8'h94;
13'd391: Q <= 8'h04;
13'd392: Q <= 8'h00;
13'd393: Q <= 8'h09;
13'd394: Q <= 8'h41;
13'd395: Q <= 8'h00;
13'd396: Q <= 8'h00;
13'd397: Q <= 8'h01;
13'd398: Q <= 8'h00;
13'd399: Q <= 8'h00;
13'd400: Q <= 8'haa;
13'd401: Q <= 8'ha3;
13'd402: Q <= 8'haa;
13'd403: Q <= 8'ha8;
13'd404: Q <= 8'h80;
13'd405: Q <= 8'h00;
13'd406: Q <= 8'h08;
13'd407: Q <= 8'h10;
13'd408: Q <= 8'h0c;
13'd409: Q <= 8'h88;
13'd410: Q <= 8'h28;
13'd411: Q <= 8'h00;
13'd412: Q <= 8'h00;
13'd413: Q <= 8'h00;
13'd414: Q <= 8'h08;
13'd415: Q <= 8'h00;
13'd416: Q <= 8'h10;
13'd417: Q <= 8'h32;
13'd418: Q <= 8'h00;
13'd419: Q <= 8'h00;
13'd420: Q <= 8'h30;
13'd421: Q <= 8'h00;
13'd422: Q <= 8'h00;
13'd423: Q <= 8'h00;
13'd424: Q <= 8'h11;
13'd425: Q <= 8'h95;
13'd426: Q <= 8'h40;
13'd427: Q <= 8'h20;
13'd428: Q <= 8'h75;
13'd429: Q <= 8'h55;
13'd430: Q <= 8'h02;
13'd431: Q <= 8'h00;
13'd432: Q <= 8'h50;
13'd433: Q <= 8'h98;
13'd434: Q <= 8'h00;
13'd435: Q <= 8'h00;
13'd436: Q <= 8'h00;
13'd437: Q <= 8'h50;
13'd438: Q <= 8'h00;
13'd439: Q <= 8'h00;
13'd440: Q <= 8'h53;
13'd441: Q <= 8'h9b;
13'd442: Q <= 8'h11;
13'd443: Q <= 8'h00;
13'd444: Q <= 8'hff;
13'd445: Q <= 8'hf0;
13'd446: Q <= 8'h51;
13'd447: Q <= 8'h04;
13'd448: Q <= 8'h80;
13'd449: Q <= 8'h00;
13'd450: Q <= 8'h10;
13'd451: Q <= 8'h10;
13'd452: Q <= 8'h80;
13'd453: Q <= 8'h00;
13'd454: Q <= 8'h00;
13'd455: Q <= 8'h1b;
13'd456: Q <= 8'hf3;
13'd457: Q <= 8'h01;
13'd458: Q <= 8'h10;
13'd459: Q <= 8'h13;
13'd460: Q <= 8'h01;
13'd461: Q <= 8'h00;
13'd462: Q <= 8'h03;
13'd463: Q <= 8'h5f;
13'd464: Q <= 8'h3e;
13'd465: Q <= 8'h08;
13'd466: Q <= 8'h00;
13'd467: Q <= 8'h00;
13'd468: Q <= 8'h02;
13'd469: Q <= 8'h00;
13'd470: Q <= 8'h04;
13'd471: Q <= 8'h3b;
13'd472: Q <= 8'hbf;
13'd473: Q <= 8'h2b;
13'd474: Q <= 8'h25;
13'd475: Q <= 8'h1d;
13'd476: Q <= 8'h1c;
13'd477: Q <= 8'h08;
13'd478: Q <= 8'h0d;
13'd479: Q <= 8'h1f;
13'd480: Q <= 8'hd8;
13'd481: Q <= 8'hd6;
13'd482: Q <= 8'hc0;
13'd483: Q <= 8'hde;
13'd484: Q <= 8'h80;
13'd485: Q <= 8'h90;
13'd486: Q <= 8'h0c;
13'd487: Q <= 8'hd8;
13'd488: Q <= 8'h00;
13'd489: Q <= 8'h40;
13'd490: Q <= 8'h00;
13'd491: Q <= 8'h50;
13'd492: Q <= 8'h00;
13'd493: Q <= 8'hd0;
13'd494: Q <= 8'h20;
13'd495: Q <= 8'h40;
13'd496: Q <= 8'hc1;
13'd497: Q <= 8'he0;
13'd498: Q <= 8'he0;
13'd499: Q <= 8'h88;
13'd500: Q <= 8'h00;
13'd501: Q <= 8'h00;
13'd502: Q <= 8'h00;
13'd503: Q <= 8'hc1;
13'd504: Q <= 8'ha0;
13'd505: Q <= 8'h40;
13'd506: Q <= 8'h00;
13'd507: Q <= 8'h02;
13'd508: Q <= 8'h00;
13'd509: Q <= 8'h00;
13'd510: Q <= 8'h00;
13'd511: Q <= 8'h00;
13'd512: Q <= 8'heb;
13'd513: Q <= 8'h0a;
13'd514: Q <= 8'h00;
13'd515: Q <= 8'h20;
13'd516: Q <= 8'hca;
13'd517: Q <= 8'h48;
13'd518: Q <= 8'h89;
13'd519: Q <= 8'hcb;
13'd520: Q <= 8'h23;
13'd521: Q <= 8'h00;
13'd522: Q <= 8'h01;
13'd523: Q <= 8'h01;
13'd524: Q <= 8'h00;
13'd525: Q <= 8'h00;
13'd526: Q <= 8'h40;
13'd527: Q <= 8'h01;
13'd528: Q <= 8'hab;
13'd529: Q <= 8'h08;
13'd530: Q <= 8'h88;
13'd531: Q <= 8'h0a;
13'd532: Q <= 8'h8a;
13'd533: Q <= 8'h00;
13'd534: Q <= 8'h0a;
13'd535: Q <= 8'h0a;
13'd536: Q <= 8'h2b;
13'd537: Q <= 8'h00;
13'd538: Q <= 8'h00;
13'd539: Q <= 8'h01;
13'd540: Q <= 8'hc1;
13'd541: Q <= 8'h00;
13'd542: Q <= 8'h00;
13'd543: Q <= 8'h02;
13'd544: Q <= 8'h00;
13'd545: Q <= 8'h00;
13'd546: Q <= 8'h00;
13'd547: Q <= 8'h00;
13'd548: Q <= 8'h98;
13'd549: Q <= 8'h05;
13'd550: Q <= 8'hc1;
13'd551: Q <= 8'h03;
13'd552: Q <= 8'h99;
13'd553: Q <= 8'h19;
13'd554: Q <= 8'h01;
13'd555: Q <= 8'h41;
13'd556: Q <= 8'hdd;
13'd557: Q <= 8'h9f;
13'd558: Q <= 8'hff;
13'd559: Q <= 8'hcf;
13'd560: Q <= 8'hda;
13'd561: Q <= 8'h00;
13'd562: Q <= 8'h80;
13'd563: Q <= 8'h00;
13'd564: Q <= 8'hba;
13'd565: Q <= 8'h0a;
13'd566: Q <= 8'h80;
13'd567: Q <= 8'h02;
13'd568: Q <= 8'h98;
13'd569: Q <= 8'h9a;
13'd570: Q <= 8'h00;
13'd571: Q <= 8'h00;
13'd572: Q <= 8'h88;
13'd573: Q <= 8'h3b;
13'd574: Q <= 8'ha8;
13'd575: Q <= 8'h1f;
13'd576: Q <= 8'hb3;
13'd577: Q <= 8'h01;
13'd578: Q <= 8'h3b;
13'd579: Q <= 8'h2b;
13'd580: Q <= 8'h28;
13'd581: Q <= 8'h01;
13'd582: Q <= 8'hab;
13'd583: Q <= 8'haf;
13'd584: Q <= 8'h08;
13'd585: Q <= 8'h02;
13'd586: Q <= 8'h0d;
13'd587: Q <= 8'h00;
13'd588: Q <= 8'h08;
13'd589: Q <= 8'h80;
13'd590: Q <= 8'h00;
13'd591: Q <= 8'h01;
13'd592: Q <= 8'h33;
13'd593: Q <= 8'h38;
13'd594: Q <= 8'h32;
13'd595: Q <= 8'ha7;
13'd596: Q <= 8'h08;
13'd597: Q <= 8'h00;
13'd598: Q <= 8'h02;
13'd599: Q <= 8'h0a;
13'd600: Q <= 8'h00;
13'd601: Q <= 8'h00;
13'd602: Q <= 8'h00;
13'd603: Q <= 8'h00;
13'd604: Q <= 8'h00;
13'd605: Q <= 8'h00;
13'd606: Q <= 8'h00;
13'd607: Q <= 8'h00;
13'd608: Q <= 8'h08;
13'd609: Q <= 8'h80;
13'd610: Q <= 8'h00;
13'd611: Q <= 8'h00;
13'd612: Q <= 8'hdd;
13'd613: Q <= 8'hc4;
13'd614: Q <= 8'h00;
13'd615: Q <= 8'hc4;
13'd616: Q <= 8'h40;
13'd617: Q <= 8'h00;
13'd618: Q <= 8'h00;
13'd619: Q <= 8'h00;
13'd620: Q <= 8'hd4;
13'd621: Q <= 8'h44;
13'd622: Q <= 8'h40;
13'd623: Q <= 8'hc8;
13'd624: Q <= 8'h00;
13'd625: Q <= 8'h00;
13'd626: Q <= 8'h80;
13'd627: Q <= 8'h00;
13'd628: Q <= 8'h00;
13'd629: Q <= 8'h00;
13'd630: Q <= 8'h44;
13'd631: Q <= 8'h40;
13'd632: Q <= 8'h00;
13'd633: Q <= 8'h00;
13'd634: Q <= 8'h00;
13'd635: Q <= 8'h00;
13'd636: Q <= 8'hc4;
13'd637: Q <= 8'hc8;
13'd638: Q <= 8'h41;
13'd639: Q <= 8'hd4;
13'd640: Q <= 8'h90;
13'd641: Q <= 8'h3d;
13'd642: Q <= 8'h18;
13'd643: Q <= 8'h05;
13'd644: Q <= 8'h20;
13'd645: Q <= 8'h11;
13'd646: Q <= 8'h84;
13'd647: Q <= 8'h80;
13'd648: Q <= 8'h11;
13'd649: Q <= 8'hc5;
13'd650: Q <= 8'hc6;
13'd651: Q <= 8'h3d;
13'd652: Q <= 8'h00;
13'd653: Q <= 8'h05;
13'd654: Q <= 8'h44;
13'd655: Q <= 8'hcf;
13'd656: Q <= 8'hba;
13'd657: Q <= 8'hbf;
13'd658: Q <= 8'h0a;
13'd659: Q <= 8'hbd;
13'd660: Q <= 8'h08;
13'd661: Q <= 8'h2b;
13'd662: Q <= 8'h81;
13'd663: Q <= 8'h03;
13'd664: Q <= 8'h40;
13'd665: Q <= 8'h4d;
13'd666: Q <= 8'h68;
13'd667: Q <= 8'h3c;
13'd668: Q <= 8'h00;
13'd669: Q <= 8'h0a;
13'd670: Q <= 8'h98;
13'd671: Q <= 8'h0b;
13'd672: Q <= 8'h00;
13'd673: Q <= 8'h44;
13'd674: Q <= 8'h00;
13'd675: Q <= 8'h00;
13'd676: Q <= 8'h00;
13'd677: Q <= 8'h50;
13'd678: Q <= 8'h00;
13'd679: Q <= 8'h00;
13'd680: Q <= 8'h44;
13'd681: Q <= 8'h57;
13'd682: Q <= 8'h00;
13'd683: Q <= 8'h10;
13'd684: Q <= 8'h04;
13'd685: Q <= 8'h55;
13'd686: Q <= 8'h00;
13'd687: Q <= 8'h08;
13'd688: Q <= 8'h40;
13'd689: Q <= 8'h44;
13'd690: Q <= 8'h00;
13'd691: Q <= 8'h00;
13'd692: Q <= 8'h00;
13'd693: Q <= 8'h00;
13'd694: Q <= 8'h00;
13'd695: Q <= 8'h00;
13'd696: Q <= 8'h44;
13'd697: Q <= 8'h55;
13'd698: Q <= 8'h00;
13'd699: Q <= 8'h00;
13'd700: Q <= 8'h55;
13'd701: Q <= 8'h55;
13'd702: Q <= 8'h00;
13'd703: Q <= 8'h00;
13'd704: Q <= 8'h10;
13'd705: Q <= 8'h11;
13'd706: Q <= 8'h00;
13'd707: Q <= 8'h30;
13'd708: Q <= 8'h55;
13'd709: Q <= 8'hf1;
13'd710: Q <= 8'h10;
13'd711: Q <= 8'h7d;
13'd712: Q <= 8'hd4;
13'd713: Q <= 8'h50;
13'd714: Q <= 8'h10;
13'd715: Q <= 8'h10;
13'd716: Q <= 8'hd5;
13'd717: Q <= 8'hd5;
13'd718: Q <= 8'h51;
13'd719: Q <= 8'hd7;
13'd720: Q <= 8'h80;
13'd721: Q <= 8'h00;
13'd722: Q <= 8'h00;
13'd723: Q <= 8'h80;
13'd724: Q <= 8'h00;
13'd725: Q <= 8'hf0;
13'd726: Q <= 8'h40;
13'd727: Q <= 8'h98;
13'd728: Q <= 8'hc0;
13'd729: Q <= 8'h00;
13'd730: Q <= 8'h00;
13'd731: Q <= 8'h41;
13'd732: Q <= 8'h40;
13'd733: Q <= 8'h90;
13'd734: Q <= 8'h00;
13'd735: Q <= 8'h10;
13'd736: Q <= 8'h2d;
13'd737: Q <= 8'h03;
13'd738: Q <= 8'h00;
13'd739: Q <= 8'h04;
13'd740: Q <= 8'h00;
13'd741: Q <= 8'h18;
13'd742: Q <= 8'h00;
13'd743: Q <= 8'h00;
13'd744: Q <= 8'h07;
13'd745: Q <= 8'h00;
13'd746: Q <= 8'h00;
13'd747: Q <= 8'h00;
13'd748: Q <= 8'h27;
13'd749: Q <= 8'h03;
13'd750: Q <= 8'h3d;
13'd751: Q <= 8'h05;
13'd752: Q <= 8'h00;
13'd753: Q <= 8'h50;
13'd754: Q <= 8'h00;
13'd755: Q <= 8'h00;
13'd756: Q <= 8'h00;
13'd757: Q <= 8'h50;
13'd758: Q <= 8'h00;
13'd759: Q <= 8'h40;
13'd760: Q <= 8'h17;
13'd761: Q <= 8'h01;
13'd762: Q <= 8'h08;
13'd763: Q <= 8'h03;
13'd764: Q <= 8'h1f;
13'd765: Q <= 8'h1b;
13'd766: Q <= 8'h01;
13'd767: Q <= 8'h01;
13'd768: Q <= 8'hd8;
13'd769: Q <= 8'h40;
13'd770: Q <= 8'h40;
13'd771: Q <= 8'h08;
13'd772: Q <= 8'h08;
13'd773: Q <= 8'h50;
13'd774: Q <= 8'h40;
13'd775: Q <= 8'hc4;
13'd776: Q <= 8'hf4;
13'd777: Q <= 8'hd1;
13'd778: Q <= 8'h00;
13'd779: Q <= 8'h51;
13'd780: Q <= 8'h00;
13'd781: Q <= 8'h00;
13'd782: Q <= 8'hc4;
13'd783: Q <= 8'h71;
13'd784: Q <= 8'hdd;
13'd785: Q <= 8'hcb;
13'd786: Q <= 8'h44;
13'd787: Q <= 8'h50;
13'd788: Q <= 8'h08;
13'd789: Q <= 8'h00;
13'd790: Q <= 8'hc1;
13'd791: Q <= 8'hc9;
13'd792: Q <= 8'hd7;
13'd793: Q <= 8'hda;
13'd794: Q <= 8'h00;
13'd795: Q <= 8'h51;
13'd796: Q <= 8'h48;
13'd797: Q <= 8'h00;
13'd798: Q <= 8'h40;
13'd799: Q <= 8'h50;
13'd800: Q <= 8'h50;
13'd801: Q <= 8'h25;
13'd802: Q <= 8'h50;
13'd803: Q <= 8'h05;
13'd804: Q <= 8'h00;
13'd805: Q <= 8'h08;
13'd806: Q <= 8'h40;
13'd807: Q <= 8'h00;
13'd808: Q <= 8'h25;
13'd809: Q <= 8'hd9;
13'd810: Q <= 8'h1a;
13'd811: Q <= 8'hb5;
13'd812: Q <= 8'hd1;
13'd813: Q <= 8'h57;
13'd814: Q <= 8'h50;
13'd815: Q <= 8'h4f;
13'd816: Q <= 8'hda;
13'd817: Q <= 8'h9b;
13'd818: Q <= 8'h80;
13'd819: Q <= 8'hb7;
13'd820: Q <= 8'ha8;
13'd821: Q <= 8'h39;
13'd822: Q <= 8'h28;
13'd823: Q <= 8'h02;
13'd824: Q <= 8'ha9;
13'd825: Q <= 8'hdb;
13'd826: Q <= 8'h00;
13'd827: Q <= 8'hfe;
13'd828: Q <= 8'h98;
13'd829: Q <= 8'h3b;
13'd830: Q <= 8'h0c;
13'd831: Q <= 8'h09;
13'd832: Q <= 8'h97;
13'd833: Q <= 8'h93;
13'd834: Q <= 8'hff;
13'd835: Q <= 8'hbf;
13'd836: Q <= 8'h02;
13'd837: Q <= 8'h82;
13'd838: Q <= 8'haf;
13'd839: Q <= 8'hf3;
13'd840: Q <= 8'h08;
13'd841: Q <= 8'h01;
13'd842: Q <= 8'h07;
13'd843: Q <= 8'h02;
13'd844: Q <= 8'h00;
13'd845: Q <= 8'h00;
13'd846: Q <= 8'h00;
13'd847: Q <= 8'h02;
13'd848: Q <= 8'h13;
13'd849: Q <= 8'h07;
13'd850: Q <= 8'h0f;
13'd851: Q <= 8'h2f;
13'd852: Q <= 8'h80;
13'd853: Q <= 8'h00;
13'd854: Q <= 8'h0b;
13'd855: Q <= 8'h06;
13'd856: Q <= 8'h00;
13'd857: Q <= 8'h00;
13'd858: Q <= 8'h24;
13'd859: Q <= 8'h29;
13'd860: Q <= 8'h00;
13'd861: Q <= 8'h08;
13'd862: Q <= 8'h04;
13'd863: Q <= 8'h00;
13'd864: Q <= 8'h04;
13'd865: Q <= 8'hca;
13'd866: Q <= 8'h5f;
13'd867: Q <= 8'h55;
13'd868: Q <= 8'h00;
13'd869: Q <= 8'h80;
13'd870: Q <= 8'h17;
13'd871: Q <= 8'h31;
13'd872: Q <= 8'h00;
13'd873: Q <= 8'hc0;
13'd874: Q <= 8'h00;
13'd875: Q <= 8'h00;
13'd876: Q <= 8'h0b;
13'd877: Q <= 8'h40;
13'd878: Q <= 8'h0b;
13'd879: Q <= 8'h02;
13'd880: Q <= 8'h02;
13'd881: Q <= 8'h00;
13'd882: Q <= 8'h10;
13'd883: Q <= 8'h10;
13'd884: Q <= 8'h00;
13'd885: Q <= 8'h00;
13'd886: Q <= 8'h09;
13'd887: Q <= 8'h50;
13'd888: Q <= 8'h00;
13'd889: Q <= 8'h00;
13'd890: Q <= 8'h44;
13'd891: Q <= 8'h40;
13'd892: Q <= 8'h02;
13'd893: Q <= 8'h80;
13'd894: Q <= 8'h13;
13'd895: Q <= 8'h00;
13'd896: Q <= 8'hcf;
13'd897: Q <= 8'h00;
13'd898: Q <= 8'h9f;
13'd899: Q <= 8'h3f;
13'd900: Q <= 8'h80;
13'd901: Q <= 8'h08;
13'd902: Q <= 8'hab;
13'd903: Q <= 8'h0b;
13'd904: Q <= 8'h88;
13'd905: Q <= 8'h40;
13'd906: Q <= 8'h08;
13'd907: Q <= 8'h1a;
13'd908: Q <= 8'h02;
13'd909: Q <= 8'h00;
13'd910: Q <= 8'h00;
13'd911: Q <= 8'h08;
13'd912: Q <= 8'h33;
13'd913: Q <= 8'h00;
13'd914: Q <= 8'h08;
13'd915: Q <= 8'h03;
13'd916: Q <= 8'h80;
13'd917: Q <= 8'h00;
13'd918: Q <= 8'h00;
13'd919: Q <= 8'h00;
13'd920: Q <= 8'h00;
13'd921: Q <= 8'h00;
13'd922: Q <= 8'h00;
13'd923: Q <= 8'h00;
13'd924: Q <= 8'h00;
13'd925: Q <= 8'h00;
13'd926: Q <= 8'h00;
13'd927: Q <= 8'h00;
13'd928: Q <= 8'hca;
13'd929: Q <= 8'h88;
13'd930: Q <= 8'h60;
13'd931: Q <= 8'hce;
13'd932: Q <= 8'h42;
13'd933: Q <= 8'h80;
13'd934: Q <= 8'h08;
13'd935: Q <= 8'h02;
13'd936: Q <= 8'h00;
13'd937: Q <= 8'h80;
13'd938: Q <= 8'h8d;
13'd939: Q <= 8'h01;
13'd940: Q <= 8'h00;
13'd941: Q <= 8'h88;
13'd942: Q <= 8'h40;
13'd943: Q <= 8'h19;
13'd944: Q <= 8'h8b;
13'd945: Q <= 8'h80;
13'd946: Q <= 8'h00;
13'd947: Q <= 8'h10;
13'd948: Q <= 8'h80;
13'd949: Q <= 8'h08;
13'd950: Q <= 8'h88;
13'd951: Q <= 8'h82;
13'd952: Q <= 8'hc3;
13'd953: Q <= 8'h42;
13'd954: Q <= 8'h20;
13'd955: Q <= 8'h00;
13'd956: Q <= 8'h90;
13'd957: Q <= 8'h00;
13'd958: Q <= 8'h09;
13'd959: Q <= 8'h01;
13'd960: Q <= 8'h8f;
13'd961: Q <= 8'h88;
13'd962: Q <= 8'hef;
13'd963: Q <= 8'h40;
13'd964: Q <= 8'h40;
13'd965: Q <= 8'h80;
13'd966: Q <= 8'h67;
13'd967: Q <= 8'h40;
13'd968: Q <= 8'h00;
13'd969: Q <= 8'h80;
13'd970: Q <= 8'h43;
13'd971: Q <= 8'h80;
13'd972: Q <= 8'h08;
13'd973: Q <= 8'h00;
13'd974: Q <= 8'h11;
13'd975: Q <= 8'h00;
13'd976: Q <= 8'h0b;
13'd977: Q <= 8'h80;
13'd978: Q <= 8'h01;
13'd979: Q <= 8'h44;
13'd980: Q <= 8'h02;
13'd981: Q <= 8'h00;
13'd982: Q <= 8'h00;
13'd983: Q <= 8'h00;
13'd984: Q <= 8'h0b;
13'd985: Q <= 8'h08;
13'd986: Q <= 8'h24;
13'd987: Q <= 8'h00;
13'd988: Q <= 8'hbb;
13'd989: Q <= 8'h48;
13'd990: Q <= 8'h0b;
13'd991: Q <= 8'h00;
13'd992: Q <= 8'h00;
13'd993: Q <= 8'h08;
13'd994: Q <= 8'h05;
13'd995: Q <= 8'h40;
13'd996: Q <= 8'h00;
13'd997: Q <= 8'h00;
13'd998: Q <= 8'h04;
13'd999: Q <= 8'h40;
13'd1000: Q <= 8'h00;
13'd1001: Q <= 8'h00;
13'd1002: Q <= 8'h00;
13'd1003: Q <= 8'h00;
13'd1004: Q <= 8'h05;
13'd1005: Q <= 8'h51;
13'd1006: Q <= 8'h4d;
13'd1007: Q <= 8'h4c;
13'd1008: Q <= 8'h10;
13'd1009: Q <= 8'h40;
13'd1010: Q <= 8'h51;
13'd1011: Q <= 8'h00;
13'd1012: Q <= 8'h00;
13'd1013: Q <= 8'h00;
13'd1014: Q <= 8'h00;
13'd1015: Q <= 8'h00;
13'd1016: Q <= 8'h41;
13'd1017: Q <= 8'h10;
13'd1018: Q <= 8'h00;
13'd1019: Q <= 8'h14;
13'd1020: Q <= 8'h55;
13'd1021: Q <= 8'h55;
13'd1022: Q <= 8'h4d;
13'd1023: Q <= 8'hdd;
13'd1024: Q <= 8'h33;
13'd1025: Q <= 8'h02;
13'd1026: Q <= 8'h23;
13'd1027: Q <= 8'h2a;
13'd1028: Q <= 8'h63;
13'd1029: Q <= 8'h00;
13'd1030: Q <= 8'h0b;
13'd1031: Q <= 8'h2a;
13'd1032: Q <= 8'h53;
13'd1033: Q <= 8'h00;
13'd1034: Q <= 8'h30;
13'd1035: Q <= 8'h20;
13'd1036: Q <= 8'h32;
13'd1037: Q <= 8'h10;
13'd1038: Q <= 8'h01;
13'd1039: Q <= 8'h22;
13'd1040: Q <= 8'h02;
13'd1041: Q <= 8'h22;
13'd1042: Q <= 8'h03;
13'd1043: Q <= 8'h22;
13'd1044: Q <= 8'h2a;
13'd1045: Q <= 8'h00;
13'd1046: Q <= 8'h0a;
13'd1047: Q <= 8'h23;
13'd1048: Q <= 8'h03;
13'd1049: Q <= 8'h20;
13'd1050: Q <= 8'h01;
13'd1051: Q <= 8'h02;
13'd1052: Q <= 8'h00;
13'd1053: Q <= 8'h00;
13'd1054: Q <= 8'h23;
13'd1055: Q <= 8'h02;
13'd1056: Q <= 8'h0c;
13'd1057: Q <= 8'h40;
13'd1058: Q <= 8'h55;
13'd1059: Q <= 8'h79;
13'd1060: Q <= 8'h09;
13'd1061: Q <= 8'h50;
13'd1062: Q <= 8'h7d;
13'd1063: Q <= 8'hfd;
13'd1064: Q <= 8'h0c;
13'd1065: Q <= 8'h08;
13'd1066: Q <= 8'h01;
13'd1067: Q <= 8'h10;
13'd1068: Q <= 8'h13;
13'd1069: Q <= 8'h81;
13'd1070: Q <= 8'h19;
13'd1071: Q <= 8'h00;
13'd1072: Q <= 8'h00;
13'd1073: Q <= 8'h30;
13'd1074: Q <= 8'h71;
13'd1075: Q <= 8'hf0;
13'd1076: Q <= 8'h10;
13'd1077: Q <= 8'h80;
13'd1078: Q <= 8'hff;
13'd1079: Q <= 8'hb0;
13'd1080: Q <= 8'h00;
13'd1081: Q <= 8'h50;
13'd1082: Q <= 8'h82;
13'd1083: Q <= 8'h8b;
13'd1084: Q <= 8'h50;
13'd1085: Q <= 8'h00;
13'd1086: Q <= 8'h00;
13'd1087: Q <= 8'h30;
13'd1088: Q <= 8'hcf;
13'd1089: Q <= 8'h0e;
13'd1090: Q <= 8'hd7;
13'd1091: Q <= 8'h10;
13'd1092: Q <= 8'hff;
13'd1093: Q <= 8'h4e;
13'd1094: Q <= 8'hde;
13'd1095: Q <= 8'h5c;
13'd1096: Q <= 8'h4f;
13'd1097: Q <= 8'hae;
13'd1098: Q <= 8'h00;
13'd1099: Q <= 8'hab;
13'd1100: Q <= 8'hef;
13'd1101: Q <= 8'h06;
13'd1102: Q <= 8'h2a;
13'd1103: Q <= 8'h0a;
13'd1104: Q <= 8'h66;
13'd1105: Q <= 8'h00;
13'd1106: Q <= 8'h98;
13'd1107: Q <= 8'h20;
13'd1108: Q <= 8'hcc;
13'd1109: Q <= 8'h04;
13'd1110: Q <= 8'h4e;
13'd1111: Q <= 8'h00;
13'd1112: Q <= 8'h2e;
13'd1113: Q <= 8'h83;
13'd1114: Q <= 8'h0a;
13'd1115: Q <= 8'h02;
13'd1116: Q <= 8'h18;
13'd1117: Q <= 8'h0a;
13'd1118: Q <= 8'h00;
13'd1119: Q <= 8'h22;
13'd1120: Q <= 8'h2b;
13'd1121: Q <= 8'hff;
13'd1122: Q <= 8'h6b;
13'd1123: Q <= 8'hc3;
13'd1124: Q <= 8'h0a;
13'd1125: Q <= 8'h6e;
13'd1126: Q <= 8'h23;
13'd1127: Q <= 8'h24;
13'd1128: Q <= 8'h02;
13'd1129: Q <= 8'hc5;
13'd1130: Q <= 8'h74;
13'd1131: Q <= 8'hc9;
13'd1132: Q <= 8'h20;
13'd1133: Q <= 8'hce;
13'd1134: Q <= 8'h60;
13'd1135: Q <= 8'h40;
13'd1136: Q <= 8'h47;
13'd1137: Q <= 8'hcf;
13'd1138: Q <= 8'h7e;
13'd1139: Q <= 8'h6d;
13'd1140: Q <= 8'h17;
13'd1141: Q <= 8'h5f;
13'd1142: Q <= 8'h28;
13'd1143: Q <= 8'h51;
13'd1144: Q <= 8'h24;
13'd1145: Q <= 8'h84;
13'd1146: Q <= 8'h02;
13'd1147: Q <= 8'h80;
13'd1148: Q <= 8'h42;
13'd1149: Q <= 8'hfc;
13'd1150: Q <= 8'h57;
13'd1151: Q <= 8'hc0;
13'd1152: Q <= 8'h45;
13'd1153: Q <= 8'h2d;
13'd1154: Q <= 8'h20;
13'd1155: Q <= 8'h27;
13'd1156: Q <= 8'h29;
13'd1157: Q <= 8'h2f;
13'd1158: Q <= 8'heb;
13'd1159: Q <= 8'h00;
13'd1160: Q <= 8'h2d;
13'd1161: Q <= 8'ha3;
13'd1162: Q <= 8'h70;
13'd1163: Q <= 8'h08;
13'd1164: Q <= 8'h3b;
13'd1165: Q <= 8'hb3;
13'd1166: Q <= 8'hf7;
13'd1167: Q <= 8'h23;
13'd1168: Q <= 8'h05;
13'd1169: Q <= 8'h05;
13'd1170: Q <= 8'h3d;
13'd1171: Q <= 8'ha6;
13'd1172: Q <= 8'h51;
13'd1173: Q <= 8'h2a;
13'd1174: Q <= 8'hf1;
13'd1175: Q <= 8'h2e;
13'd1176: Q <= 8'h4d;
13'd1177: Q <= 8'h02;
13'd1178: Q <= 8'hc2;
13'd1179: Q <= 8'h04;
13'd1180: Q <= 8'h5d;
13'd1181: Q <= 8'h31;
13'd1182: Q <= 8'h0c;
13'd1183: Q <= 8'h4f;
13'd1184: Q <= 8'hdf;
13'd1185: Q <= 8'h32;
13'd1186: Q <= 8'hbd;
13'd1187: Q <= 8'h35;
13'd1188: Q <= 8'h00;
13'd1189: Q <= 8'h00;
13'd1190: Q <= 8'h09;
13'd1191: Q <= 8'h0c;
13'd1192: Q <= 8'h05;
13'd1193: Q <= 8'h01;
13'd1194: Q <= 8'h00;
13'd1195: Q <= 8'h00;
13'd1196: Q <= 8'h00;
13'd1197: Q <= 8'h00;
13'd1198: Q <= 8'h04;
13'd1199: Q <= 8'h04;
13'd1200: Q <= 8'hef;
13'd1201: Q <= 8'hc4;
13'd1202: Q <= 8'h8a;
13'd1203: Q <= 8'h08;
13'd1204: Q <= 8'h00;
13'd1205: Q <= 8'h00;
13'd1206: Q <= 8'h08;
13'd1207: Q <= 8'h00;
13'd1208: Q <= 8'h89;
13'd1209: Q <= 8'h00;
13'd1210: Q <= 8'h80;
13'd1211: Q <= 8'h02;
13'd1212: Q <= 8'h00;
13'd1213: Q <= 8'h00;
13'd1214: Q <= 8'h00;
13'd1215: Q <= 8'h00;
13'd1216: Q <= 8'hca;
13'd1217: Q <= 8'hc8;
13'd1218: Q <= 8'h44;
13'd1219: Q <= 8'h00;
13'd1220: Q <= 8'h80;
13'd1221: Q <= 8'h90;
13'd1222: Q <= 8'h84;
13'd1223: Q <= 8'h18;
13'd1224: Q <= 8'h08;
13'd1225: Q <= 8'h08;
13'd1226: Q <= 8'h00;
13'd1227: Q <= 8'h10;
13'd1228: Q <= 8'h40;
13'd1229: Q <= 8'h00;
13'd1230: Q <= 8'h06;
13'd1231: Q <= 8'h04;
13'd1232: Q <= 8'hca;
13'd1233: Q <= 8'hc0;
13'd1234: Q <= 8'h08;
13'd1235: Q <= 8'h01;
13'd1236: Q <= 8'h84;
13'd1237: Q <= 8'h80;
13'd1238: Q <= 8'h00;
13'd1239: Q <= 8'h00;
13'd1240: Q <= 8'hba;
13'd1241: Q <= 8'ha0;
13'd1242: Q <= 8'h40;
13'd1243: Q <= 8'h04;
13'd1244: Q <= 8'hc0;
13'd1245: Q <= 8'h72;
13'd1246: Q <= 8'h00;
13'd1247: Q <= 8'h00;
13'd1248: Q <= 8'h00;
13'd1249: Q <= 8'h10;
13'd1250: Q <= 8'h86;
13'd1251: Q <= 8'h04;
13'd1252: Q <= 8'h6d;
13'd1253: Q <= 8'h11;
13'd1254: Q <= 8'hff;
13'd1255: Q <= 8'h06;
13'd1256: Q <= 8'h22;
13'd1257: Q <= 8'hd2;
13'd1258: Q <= 8'h3f;
13'd1259: Q <= 8'h0e;
13'd1260: Q <= 8'h83;
13'd1261: Q <= 8'h52;
13'd1262: Q <= 8'hbf;
13'd1263: Q <= 8'h00;
13'd1264: Q <= 8'h01;
13'd1265: Q <= 8'h99;
13'd1266: Q <= 8'h7b;
13'd1267: Q <= 8'ha7;
13'd1268: Q <= 8'h02;
13'd1269: Q <= 8'h32;
13'd1270: Q <= 8'h3f;
13'd1271: Q <= 8'h84;
13'd1272: Q <= 8'h00;
13'd1273: Q <= 8'hc7;
13'd1274: Q <= 8'h73;
13'd1275: Q <= 8'h81;
13'd1276: Q <= 8'h10;
13'd1277: Q <= 8'hdf;
13'd1278: Q <= 8'h33;
13'd1279: Q <= 8'hd0;
13'd1280: Q <= 8'h5c;
13'd1281: Q <= 8'h50;
13'd1282: Q <= 8'h15;
13'd1283: Q <= 8'h31;
13'd1284: Q <= 8'h12;
13'd1285: Q <= 8'h00;
13'd1286: Q <= 8'h1d;
13'd1287: Q <= 8'hd1;
13'd1288: Q <= 8'h10;
13'd1289: Q <= 8'h82;
13'd1290: Q <= 8'h01;
13'd1291: Q <= 8'h01;
13'd1292: Q <= 8'h01;
13'd1293: Q <= 8'h00;
13'd1294: Q <= 8'h51;
13'd1295: Q <= 8'h51;
13'd1296: Q <= 8'h24;
13'd1297: Q <= 8'hda;
13'd1298: Q <= 8'h90;
13'd1299: Q <= 8'hf1;
13'd1300: Q <= 8'h02;
13'd1301: Q <= 8'h80;
13'd1302: Q <= 8'h90;
13'd1303: Q <= 8'hb1;
13'd1304: Q <= 8'h20;
13'd1305: Q <= 8'h38;
13'd1306: Q <= 8'h80;
13'd1307: Q <= 8'h29;
13'd1308: Q <= 8'h4c;
13'd1309: Q <= 8'h03;
13'd1310: Q <= 8'h20;
13'd1311: Q <= 8'h1b;
13'd1312: Q <= 8'h7f;
13'd1313: Q <= 8'h1d;
13'd1314: Q <= 8'h14;
13'd1315: Q <= 8'h1f;
13'd1316: Q <= 8'h75;
13'd1317: Q <= 8'h0d;
13'd1318: Q <= 8'h99;
13'd1319: Q <= 8'hff;
13'd1320: Q <= 8'hfd;
13'd1321: Q <= 8'hdf;
13'd1322: Q <= 8'h38;
13'd1323: Q <= 8'h53;
13'd1324: Q <= 8'h11;
13'd1325: Q <= 8'h11;
13'd1326: Q <= 8'h80;
13'd1327: Q <= 8'h79;
13'd1328: Q <= 8'hdc;
13'd1329: Q <= 8'h38;
13'd1330: Q <= 8'h10;
13'd1331: Q <= 8'h0b;
13'd1332: Q <= 8'h04;
13'd1333: Q <= 8'h08;
13'd1334: Q <= 8'h90;
13'd1335: Q <= 8'hfc;
13'd1336: Q <= 8'hcc;
13'd1337: Q <= 8'h08;
13'd1338: Q <= 8'h88;
13'd1339: Q <= 8'h08;
13'd1340: Q <= 8'h04;
13'd1341: Q <= 8'h00;
13'd1342: Q <= 8'h10;
13'd1343: Q <= 8'h3e;
13'd1344: Q <= 8'h8c;
13'd1345: Q <= 8'h0c;
13'd1346: Q <= 8'h80;
13'd1347: Q <= 8'h1c;
13'd1348: Q <= 8'hcc;
13'd1349: Q <= 8'h19;
13'd1350: Q <= 8'hdd;
13'd1351: Q <= 8'hbf;
13'd1352: Q <= 8'hbe;
13'd1353: Q <= 8'h5f;
13'd1354: Q <= 8'h1a;
13'd1355: Q <= 8'h62;
13'd1356: Q <= 8'h9f;
13'd1357: Q <= 8'h33;
13'd1358: Q <= 8'h9f;
13'd1359: Q <= 8'hae;
13'd1360: Q <= 8'h00;
13'd1361: Q <= 8'h41;
13'd1362: Q <= 8'h40;
13'd1363: Q <= 8'h21;
13'd1364: Q <= 8'h50;
13'd1365: Q <= 8'h80;
13'd1366: Q <= 8'h40;
13'd1367: Q <= 8'h14;
13'd1368: Q <= 8'h3f;
13'd1369: Q <= 8'h0f;
13'd1370: Q <= 8'h04;
13'd1371: Q <= 8'haa;
13'd1372: Q <= 8'h8c;
13'd1373: Q <= 8'h09;
13'd1374: Q <= 8'h1c;
13'd1375: Q <= 8'h3f;
13'd1376: Q <= 8'h43;
13'd1377: Q <= 8'h02;
13'd1378: Q <= 8'haf;
13'd1379: Q <= 8'h0e;
13'd1380: Q <= 8'hff;
13'd1381: Q <= 8'h22;
13'd1382: Q <= 8'h5f;
13'd1383: Q <= 8'h62;
13'd1384: Q <= 8'h08;
13'd1385: Q <= 8'h00;
13'd1386: Q <= 8'h00;
13'd1387: Q <= 8'h60;
13'd1388: Q <= 8'h37;
13'd1389: Q <= 8'h0a;
13'd1390: Q <= 8'hfe;
13'd1391: Q <= 8'h2e;
13'd1392: Q <= 8'h82;
13'd1393: Q <= 8'h20;
13'd1394: Q <= 8'h86;
13'd1395: Q <= 8'ha8;
13'd1396: Q <= 8'h44;
13'd1397: Q <= 8'h88;
13'd1398: Q <= 8'h2a;
13'd1399: Q <= 8'h00;
13'd1400: Q <= 8'h00;
13'd1401: Q <= 8'h00;
13'd1402: Q <= 8'h02;
13'd1403: Q <= 8'ha8;
13'd1404: Q <= 8'h44;
13'd1405: Q <= 8'h61;
13'd1406: Q <= 8'h44;
13'd1407: Q <= 8'h00;
13'd1408: Q <= 8'hf2;
13'd1409: Q <= 8'h60;
13'd1410: Q <= 8'h00;
13'd1411: Q <= 8'h00;
13'd1412: Q <= 8'h40;
13'd1413: Q <= 8'h00;
13'd1414: Q <= 8'h40;
13'd1415: Q <= 8'ha2;
13'd1416: Q <= 8'h08;
13'd1417: Q <= 8'h80;
13'd1418: Q <= 8'h00;
13'd1419: Q <= 8'h01;
13'd1420: Q <= 8'h00;
13'd1421: Q <= 8'h00;
13'd1422: Q <= 8'h00;
13'd1423: Q <= 8'h04;
13'd1424: Q <= 8'heb;
13'd1425: Q <= 8'hc2;
13'd1426: Q <= 8'h0a;
13'd1427: Q <= 8'h80;
13'd1428: Q <= 8'h8a;
13'd1429: Q <= 8'h00;
13'd1430: Q <= 8'h88;
13'd1431: Q <= 8'haa;
13'd1432: Q <= 8'hbb;
13'd1433: Q <= 8'ha3;
13'd1434: Q <= 8'h02;
13'd1435: Q <= 8'h10;
13'd1436: Q <= 8'h34;
13'd1437: Q <= 8'h00;
13'd1438: Q <= 8'h14;
13'd1439: Q <= 8'h02;
13'd1440: Q <= 8'hce;
13'd1441: Q <= 8'h18;
13'd1442: Q <= 8'h1c;
13'd1443: Q <= 8'h00;
13'd1444: Q <= 8'h48;
13'd1445: Q <= 8'hd0;
13'd1446: Q <= 8'h00;
13'd1447: Q <= 8'h08;
13'd1448: Q <= 8'h00;
13'd1449: Q <= 8'h80;
13'd1450: Q <= 8'h00;
13'd1451: Q <= 8'h00;
13'd1452: Q <= 8'hc8;
13'd1453: Q <= 8'h00;
13'd1454: Q <= 8'h58;
13'd1455: Q <= 8'h00;
13'd1456: Q <= 8'h02;
13'd1457: Q <= 8'h0a;
13'd1458: Q <= 8'h11;
13'd1459: Q <= 8'h00;
13'd1460: Q <= 8'h88;
13'd1461: Q <= 8'h08;
13'd1462: Q <= 8'h00;
13'd1463: Q <= 8'h00;
13'd1464: Q <= 8'h26;
13'd1465: Q <= 8'h20;
13'd1466: Q <= 8'h00;
13'd1467: Q <= 8'h00;
13'd1468: Q <= 8'hfe;
13'd1469: Q <= 8'hbe;
13'd1470: Q <= 8'h00;
13'd1471: Q <= 8'h02;
13'd1472: Q <= 8'h84;
13'd1473: Q <= 8'h70;
13'd1474: Q <= 8'h08;
13'd1475: Q <= 8'h51;
13'd1476: Q <= 8'hc1;
13'd1477: Q <= 8'h00;
13'd1478: Q <= 8'h19;
13'd1479: Q <= 8'h51;
13'd1480: Q <= 8'h28;
13'd1481: Q <= 8'h90;
13'd1482: Q <= 8'h00;
13'd1483: Q <= 8'h40;
13'd1484: Q <= 8'h93;
13'd1485: Q <= 8'h10;
13'd1486: Q <= 8'h11;
13'd1487: Q <= 8'h10;
13'd1488: Q <= 8'h10;
13'd1489: Q <= 8'h30;
13'd1490: Q <= 8'h40;
13'd1491: Q <= 8'h30;
13'd1492: Q <= 8'h00;
13'd1493: Q <= 8'he0;
13'd1494: Q <= 8'h01;
13'd1495: Q <= 8'h98;
13'd1496: Q <= 8'h08;
13'd1497: Q <= 8'h40;
13'd1498: Q <= 8'h80;
13'd1499: Q <= 8'h02;
13'd1500: Q <= 8'h41;
13'd1501: Q <= 8'h42;
13'd1502: Q <= 8'h08;
13'd1503: Q <= 8'h08;
13'd1504: Q <= 8'hc0;
13'd1505: Q <= 8'hd8;
13'd1506: Q <= 8'h80;
13'd1507: Q <= 8'hd4;
13'd1508: Q <= 8'h0c;
13'd1509: Q <= 8'hd0;
13'd1510: Q <= 8'h00;
13'd1511: Q <= 8'h08;
13'd1512: Q <= 8'h40;
13'd1513: Q <= 8'hdd;
13'd1514: Q <= 8'h00;
13'd1515: Q <= 8'h44;
13'd1516: Q <= 8'h08;
13'd1517: Q <= 8'he1;
13'd1518: Q <= 8'h04;
13'd1519: Q <= 8'h0e;
13'd1520: Q <= 8'hc0;
13'd1521: Q <= 8'hc0;
13'd1522: Q <= 8'hc0;
13'd1523: Q <= 8'hd8;
13'd1524: Q <= 8'h00;
13'd1525: Q <= 8'h40;
13'd1526: Q <= 8'h00;
13'd1527: Q <= 8'h80;
13'd1528: Q <= 8'h40;
13'd1529: Q <= 8'hc4;
13'd1530: Q <= 8'h00;
13'd1531: Q <= 8'h44;
13'd1532: Q <= 8'h00;
13'd1533: Q <= 8'h40;
13'd1534: Q <= 8'h00;
13'd1535: Q <= 8'h00;
13'd1536: Q <= 8'h08;
13'd1537: Q <= 8'h08;
13'd1538: Q <= 8'h80;
13'd1539: Q <= 8'h12;
13'd1540: Q <= 8'h0a;
13'd1541: Q <= 8'h00;
13'd1542: Q <= 8'h13;
13'd1543: Q <= 8'h19;
13'd1544: Q <= 8'h9f;
13'd1545: Q <= 8'h07;
13'd1546: Q <= 8'h81;
13'd1547: Q <= 8'h0b;
13'd1548: Q <= 8'h80;
13'd1549: Q <= 8'h05;
13'd1550: Q <= 8'h13;
13'd1551: Q <= 8'h15;
13'd1552: Q <= 8'h29;
13'd1553: Q <= 8'h00;
13'd1554: Q <= 8'h28;
13'd1555: Q <= 8'hb8;
13'd1556: Q <= 8'h03;
13'd1557: Q <= 8'h00;
13'd1558: Q <= 8'h08;
13'd1559: Q <= 8'h3b;
13'd1560: Q <= 8'h9b;
13'd1561: Q <= 8'h3b;
13'd1562: Q <= 8'h18;
13'd1563: Q <= 8'hcb;
13'd1564: Q <= 8'h0d;
13'd1565: Q <= 8'h00;
13'd1566: Q <= 8'h11;
13'd1567: Q <= 8'h19;
13'd1568: Q <= 8'h00;
13'd1569: Q <= 8'h1d;
13'd1570: Q <= 8'h10;
13'd1571: Q <= 8'h55;
13'd1572: Q <= 8'h00;
13'd1573: Q <= 8'h10;
13'd1574: Q <= 8'h0c;
13'd1575: Q <= 8'h8a;
13'd1576: Q <= 8'h75;
13'd1577: Q <= 8'h19;
13'd1578: Q <= 8'h1d;
13'd1579: Q <= 8'h11;
13'd1580: Q <= 8'h11;
13'd1581: Q <= 8'h15;
13'd1582: Q <= 8'h08;
13'd1583: Q <= 8'h1d;
13'd1584: Q <= 8'hb2;
13'd1585: Q <= 8'he9;
13'd1586: Q <= 8'h28;
13'd1587: Q <= 8'hf9;
13'd1588: Q <= 8'h02;
13'd1589: Q <= 8'h91;
13'd1590: Q <= 8'h38;
13'd1591: Q <= 8'h20;
13'd1592: Q <= 8'hf2;
13'd1593: Q <= 8'hbf;
13'd1594: Q <= 8'h2b;
13'd1595: Q <= 8'h2a;
13'd1596: Q <= 8'ha4;
13'd1597: Q <= 8'hb9;
13'd1598: Q <= 8'h08;
13'd1599: Q <= 8'h28;
13'd1600: Q <= 8'h11;
13'd1601: Q <= 8'h10;
13'd1602: Q <= 8'h04;
13'd1603: Q <= 8'h2c;
13'd1604: Q <= 8'h60;
13'd1605: Q <= 8'h8c;
13'd1606: Q <= 8'h0b;
13'd1607: Q <= 8'h35;
13'd1608: Q <= 8'h7b;
13'd1609: Q <= 8'h7d;
13'd1610: Q <= 8'h91;
13'd1611: Q <= 8'h13;
13'd1612: Q <= 8'h01;
13'd1613: Q <= 8'h04;
13'd1614: Q <= 8'h43;
13'd1615: Q <= 8'h07;
13'd1616: Q <= 8'heb;
13'd1617: Q <= 8'h94;
13'd1618: Q <= 8'h1b;
13'd1619: Q <= 8'h44;
13'd1620: Q <= 8'hee;
13'd1621: Q <= 8'heb;
13'd1622: Q <= 8'h13;
13'd1623: Q <= 8'h6f;
13'd1624: Q <= 8'h36;
13'd1625: Q <= 8'h45;
13'd1626: Q <= 8'h10;
13'd1627: Q <= 8'h80;
13'd1628: Q <= 8'h10;
13'd1629: Q <= 8'h04;
13'd1630: Q <= 8'h04;
13'd1631: Q <= 8'h00;
13'd1632: Q <= 8'hab;
13'd1633: Q <= 8'h28;
13'd1634: Q <= 8'h8b;
13'd1635: Q <= 8'h04;
13'd1636: Q <= 8'h01;
13'd1637: Q <= 8'h00;
13'd1638: Q <= 8'h01;
13'd1639: Q <= 8'h00;
13'd1640: Q <= 8'h00;
13'd1641: Q <= 8'h00;
13'd1642: Q <= 8'h00;
13'd1643: Q <= 8'h00;
13'd1644: Q <= 8'h00;
13'd1645: Q <= 8'h00;
13'd1646: Q <= 8'h01;
13'd1647: Q <= 8'h04;
13'd1648: Q <= 8'h26;
13'd1649: Q <= 8'h42;
13'd1650: Q <= 8'h02;
13'd1651: Q <= 8'h00;
13'd1652: Q <= 8'h20;
13'd1653: Q <= 8'h00;
13'd1654: Q <= 8'h00;
13'd1655: Q <= 8'h00;
13'd1656: Q <= 8'h63;
13'd1657: Q <= 8'h62;
13'd1658: Q <= 8'h03;
13'd1659: Q <= 8'h00;
13'd1660: Q <= 8'hab;
13'd1661: Q <= 8'h40;
13'd1662: Q <= 8'h43;
13'd1663: Q <= 8'h10;
13'd1664: Q <= 8'hcf;
13'd1665: Q <= 8'h40;
13'd1666: Q <= 8'hff;
13'd1667: Q <= 8'he9;
13'd1668: Q <= 8'hef;
13'd1669: Q <= 8'h12;
13'd1670: Q <= 8'hdf;
13'd1671: Q <= 8'h60;
13'd1672: Q <= 8'hcb;
13'd1673: Q <= 8'h02;
13'd1674: Q <= 8'h88;
13'd1675: Q <= 8'h80;
13'd1676: Q <= 8'h0b;
13'd1677: Q <= 8'h28;
13'd1678: Q <= 8'h12;
13'd1679: Q <= 8'h00;
13'd1680: Q <= 8'hcc;
13'd1681: Q <= 8'hc0;
13'd1682: Q <= 8'hde;
13'd1683: Q <= 8'hd0;
13'd1684: Q <= 8'h06;
13'd1685: Q <= 8'h02;
13'd1686: Q <= 8'h47;
13'd1687: Q <= 8'h48;
13'd1688: Q <= 8'h50;
13'd1689: Q <= 8'hc0;
13'd1690: Q <= 8'h51;
13'd1691: Q <= 8'hd0;
13'd1692: Q <= 8'h22;
13'd1693: Q <= 8'h00;
13'd1694: Q <= 8'h44;
13'd1695: Q <= 8'h00;
13'd1696: Q <= 8'he0;
13'd1697: Q <= 8'hd0;
13'd1698: Q <= 8'h41;
13'd1699: Q <= 8'hd1;
13'd1700: Q <= 8'h08;
13'd1701: Q <= 8'h48;
13'd1702: Q <= 8'h49;
13'd1703: Q <= 8'h11;
13'd1704: Q <= 8'he0;
13'd1705: Q <= 8'h94;
13'd1706: Q <= 8'h00;
13'd1707: Q <= 8'he0;
13'd1708: Q <= 8'h02;
13'd1709: Q <= 8'h10;
13'd1710: Q <= 8'h05;
13'd1711: Q <= 8'h18;
13'd1712: Q <= 8'h8e;
13'd1713: Q <= 8'ha0;
13'd1714: Q <= 8'h03;
13'd1715: Q <= 8'h50;
13'd1716: Q <= 8'h00;
13'd1717: Q <= 8'h10;
13'd1718: Q <= 8'h00;
13'd1719: Q <= 8'h32;
13'd1720: Q <= 8'h80;
13'd1721: Q <= 8'hb2;
13'd1722: Q <= 8'h02;
13'd1723: Q <= 8'h00;
13'd1724: Q <= 8'hc0;
13'd1725: Q <= 8'h50;
13'd1726: Q <= 8'h00;
13'd1727: Q <= 8'h10;
13'd1728: Q <= 8'hff;
13'd1729: Q <= 8'h28;
13'd1730: Q <= 8'hfe;
13'd1731: Q <= 8'h1c;
13'd1732: Q <= 8'h3e;
13'd1733: Q <= 8'h38;
13'd1734: Q <= 8'h3f;
13'd1735: Q <= 8'h0a;
13'd1736: Q <= 8'hf3;
13'd1737: Q <= 8'h7c;
13'd1738: Q <= 8'h48;
13'd1739: Q <= 8'h14;
13'd1740: Q <= 8'hb1;
13'd1741: Q <= 8'h55;
13'd1742: Q <= 8'h00;
13'd1743: Q <= 8'h00;
13'd1744: Q <= 8'h0f;
13'd1745: Q <= 8'h00;
13'd1746: Q <= 8'hfb;
13'd1747: Q <= 8'h1e;
13'd1748: Q <= 8'h43;
13'd1749: Q <= 8'h3f;
13'd1750: Q <= 8'h0f;
13'd1751: Q <= 8'h2e;
13'd1752: Q <= 8'h7b;
13'd1753: Q <= 8'h5b;
13'd1754: Q <= 8'h5b;
13'd1755: Q <= 8'h04;
13'd1756: Q <= 8'h7e;
13'd1757: Q <= 8'h50;
13'd1758: Q <= 8'he3;
13'd1759: Q <= 8'h22;
13'd1760: Q <= 8'h08;
13'd1761: Q <= 8'h02;
13'd1762: Q <= 8'h00;
13'd1763: Q <= 8'h02;
13'd1764: Q <= 8'h10;
13'd1765: Q <= 8'h00;
13'd1766: Q <= 8'h55;
13'd1767: Q <= 8'h1c;
13'd1768: Q <= 8'h8f;
13'd1769: Q <= 8'h55;
13'd1770: Q <= 8'hd8;
13'd1771: Q <= 8'h54;
13'd1772: Q <= 8'h54;
13'd1773: Q <= 8'h05;
13'd1774: Q <= 8'hd0;
13'd1775: Q <= 8'h7b;
13'd1776: Q <= 8'h04;
13'd1777: Q <= 8'h00;
13'd1778: Q <= 8'h4a;
13'd1779: Q <= 8'h00;
13'd1780: Q <= 8'h44;
13'd1781: Q <= 8'h00;
13'd1782: Q <= 8'h02;
13'd1783: Q <= 8'h7c;
13'd1784: Q <= 8'h5f;
13'd1785: Q <= 8'h2d;
13'd1786: Q <= 8'h0e;
13'd1787: Q <= 8'h0d;
13'd1788: Q <= 8'h54;
13'd1789: Q <= 8'h21;
13'd1790: Q <= 8'he4;
13'd1791: Q <= 8'h3f;
13'd1792: Q <= 8'h23;
13'd1793: Q <= 8'hd2;
13'd1794: Q <= 8'hb7;
13'd1795: Q <= 8'h31;
13'd1796: Q <= 8'h03;
13'd1797: Q <= 8'hff;
13'd1798: Q <= 8'hff;
13'd1799: Q <= 8'h07;
13'd1800: Q <= 8'h22;
13'd1801: Q <= 8'he6;
13'd1802: Q <= 8'h6c;
13'd1803: Q <= 8'h50;
13'd1804: Q <= 8'h26;
13'd1805: Q <= 8'hf1;
13'd1806: Q <= 8'h00;
13'd1807: Q <= 8'h40;
13'd1808: Q <= 8'h23;
13'd1809: Q <= 8'h22;
13'd1810: Q <= 8'hf3;
13'd1811: Q <= 8'h24;
13'd1812: Q <= 8'h43;
13'd1813: Q <= 8'hff;
13'd1814: Q <= 8'h5f;
13'd1815: Q <= 8'h56;
13'd1816: Q <= 8'h50;
13'd1817: Q <= 8'h44;
13'd1818: Q <= 8'haa;
13'd1819: Q <= 8'h52;
13'd1820: Q <= 8'h56;
13'd1821: Q <= 8'hf3;
13'd1822: Q <= 8'hf6;
13'd1823: Q <= 8'h75;
13'd1824: Q <= 8'hf2;
13'd1825: Q <= 8'h90;
13'd1826: Q <= 8'h00;
13'd1827: Q <= 8'h11;
13'd1828: Q <= 8'h00;
13'd1829: Q <= 8'h80;
13'd1830: Q <= 8'h00;
13'd1831: Q <= 8'h8e;
13'd1832: Q <= 8'h91;
13'd1833: Q <= 8'h40;
13'd1834: Q <= 8'h00;
13'd1835: Q <= 8'h00;
13'd1836: Q <= 8'h15;
13'd1837: Q <= 8'h50;
13'd1838: Q <= 8'h2d;
13'd1839: Q <= 8'h67;
13'd1840: Q <= 8'h11;
13'd1841: Q <= 8'h40;
13'd1842: Q <= 8'h41;
13'd1843: Q <= 8'h45;
13'd1844: Q <= 8'h10;
13'd1845: Q <= 8'h00;
13'd1846: Q <= 8'h00;
13'd1847: Q <= 8'h50;
13'd1848: Q <= 8'h51;
13'd1849: Q <= 8'h10;
13'd1850: Q <= 8'h00;
13'd1851: Q <= 8'h10;
13'd1852: Q <= 8'h73;
13'd1853: Q <= 8'h11;
13'd1854: Q <= 8'h44;
13'd1855: Q <= 8'h57;
13'd1856: Q <= 8'h00;
13'd1857: Q <= 8'h00;
13'd1858: Q <= 8'hb8;
13'd1859: Q <= 8'hb5;
13'd1860: Q <= 8'hdd;
13'd1861: Q <= 8'h01;
13'd1862: Q <= 8'hbf;
13'd1863: Q <= 8'hbf;
13'd1864: Q <= 8'h30;
13'd1865: Q <= 8'h00;
13'd1866: Q <= 8'h99;
13'd1867: Q <= 8'h00;
13'd1868: Q <= 8'h39;
13'd1869: Q <= 8'h15;
13'd1870: Q <= 8'hff;
13'd1871: Q <= 8'hff;
13'd1872: Q <= 8'h00;
13'd1873: Q <= 8'h00;
13'd1874: Q <= 8'h88;
13'd1875: Q <= 8'h10;
13'd1876: Q <= 8'h0a;
13'd1877: Q <= 8'h00;
13'd1878: Q <= 8'h9a;
13'd1879: Q <= 8'h02;
13'd1880: Q <= 8'ha0;
13'd1881: Q <= 8'h00;
13'd1882: Q <= 8'h28;
13'd1883: Q <= 8'h48;
13'd1884: Q <= 8'hf0;
13'd1885: Q <= 8'h00;
13'd1886: Q <= 8'hba;
13'd1887: Q <= 8'hb8;
13'd1888: Q <= 8'h13;
13'd1889: Q <= 8'h3e;
13'd1890: Q <= 8'h68;
13'd1891: Q <= 8'h2e;
13'd1892: Q <= 8'h11;
13'd1893: Q <= 8'h6f;
13'd1894: Q <= 8'h88;
13'd1895: Q <= 8'h24;
13'd1896: Q <= 8'h51;
13'd1897: Q <= 8'h6b;
13'd1898: Q <= 8'h7f;
13'd1899: Q <= 8'h22;
13'd1900: Q <= 8'h7d;
13'd1901: Q <= 8'h97;
13'd1902: Q <= 8'h3d;
13'd1903: Q <= 8'h00;
13'd1904: Q <= 8'h10;
13'd1905: Q <= 8'h76;
13'd1906: Q <= 8'h06;
13'd1907: Q <= 8'h74;
13'd1908: Q <= 8'h69;
13'd1909: Q <= 8'hed;
13'd1910: Q <= 8'h6c;
13'd1911: Q <= 8'h45;
13'd1912: Q <= 8'h20;
13'd1913: Q <= 8'h70;
13'd1914: Q <= 8'h6a;
13'd1915: Q <= 8'h76;
13'd1916: Q <= 8'hae;
13'd1917: Q <= 8'haf;
13'd1918: Q <= 8'hb8;
13'd1919: Q <= 8'h00;
13'd1920: Q <= 8'hd4;
13'd1921: Q <= 8'h44;
13'd1922: Q <= 8'h00;
13'd1923: Q <= 8'h40;
13'd1924: Q <= 8'h80;
13'd1925: Q <= 8'h85;
13'd1926: Q <= 8'h00;
13'd1927: Q <= 8'h88;
13'd1928: Q <= 8'h10;
13'd1929: Q <= 8'h51;
13'd1930: Q <= 8'h40;
13'd1931: Q <= 8'h51;
13'd1932: Q <= 8'h40;
13'd1933: Q <= 8'h04;
13'd1934: Q <= 8'h85;
13'd1935: Q <= 8'h40;
13'd1936: Q <= 8'hd4;
13'd1937: Q <= 8'h4c;
13'd1938: Q <= 8'h4c;
13'd1939: Q <= 8'h54;
13'd1940: Q <= 8'h80;
13'd1941: Q <= 8'h88;
13'd1942: Q <= 8'h40;
13'd1943: Q <= 8'hcc;
13'd1944: Q <= 8'hd4;
13'd1945: Q <= 8'hf4;
13'd1946: Q <= 8'hd4;
13'd1947: Q <= 8'h50;
13'd1948: Q <= 8'h80;
13'd1949: Q <= 8'h00;
13'd1950: Q <= 8'h40;
13'd1951: Q <= 8'h40;
13'd1952: Q <= 8'h8c;
13'd1953: Q <= 8'h00;
13'd1954: Q <= 8'h04;
13'd1955: Q <= 8'h05;
13'd1956: Q <= 8'hf9;
13'd1957: Q <= 8'h04;
13'd1958: Q <= 8'hc7;
13'd1959: Q <= 8'h7c;
13'd1960: Q <= 8'h5f;
13'd1961: Q <= 8'h8e;
13'd1962: Q <= 8'hd0;
13'd1963: Q <= 8'h47;
13'd1964: Q <= 8'h04;
13'd1965: Q <= 8'h9d;
13'd1966: Q <= 8'h5d;
13'd1967: Q <= 8'hde;
13'd1968: Q <= 8'h44;
13'd1969: Q <= 8'h30;
13'd1970: Q <= 8'h00;
13'd1971: Q <= 8'h04;
13'd1972: Q <= 8'h45;
13'd1973: Q <= 8'h00;
13'd1974: Q <= 8'h00;
13'd1975: Q <= 8'h50;
13'd1976: Q <= 8'h7d;
13'd1977: Q <= 8'hbe;
13'd1978: Q <= 8'h08;
13'd1979: Q <= 8'h4e;
13'd1980: Q <= 8'h4c;
13'd1981: Q <= 8'h08;
13'd1982: Q <= 8'h4c;
13'd1983: Q <= 8'h2e;
13'd1984: Q <= 8'hf9;
13'd1985: Q <= 8'h10;
13'd1986: Q <= 8'h88;
13'd1987: Q <= 8'h01;
13'd1988: Q <= 8'h10;
13'd1989: Q <= 8'h11;
13'd1990: Q <= 8'h00;
13'd1991: Q <= 8'hfc;
13'd1992: Q <= 8'h55;
13'd1993: Q <= 8'h59;
13'd1994: Q <= 8'h4c;
13'd1995: Q <= 8'h11;
13'd1996: Q <= 8'h5c;
13'd1997: Q <= 8'h11;
13'd1998: Q <= 8'h0c;
13'd1999: Q <= 8'h0a;
13'd2000: Q <= 8'hbd;
13'd2001: Q <= 8'h8d;
13'd2002: Q <= 8'hca;
13'd2003: Q <= 8'h83;
13'd2004: Q <= 8'he0;
13'd2005: Q <= 8'h82;
13'd2006: Q <= 8'h81;
13'd2007: Q <= 8'h9a;
13'd2008: Q <= 8'hdb;
13'd2009: Q <= 8'h31;
13'd2010: Q <= 8'h98;
13'd2011: Q <= 8'h08;
13'd2012: Q <= 8'h71;
13'd2013: Q <= 8'h04;
13'd2014: Q <= 8'h00;
13'd2015: Q <= 8'h0e;
13'd2016: Q <= 8'ha3;
13'd2017: Q <= 8'hbf;
13'd2018: Q <= 8'h23;
13'd2019: Q <= 8'h33;
13'd2020: Q <= 8'h0a;
13'd2021: Q <= 8'ha3;
13'd2022: Q <= 8'h13;
13'd2023: Q <= 8'hca;
13'd2024: Q <= 8'h00;
13'd2025: Q <= 8'h40;
13'd2026: Q <= 8'h19;
13'd2027: Q <= 8'h60;
13'd2028: Q <= 8'h88;
13'd2029: Q <= 8'hb2;
13'd2030: Q <= 8'h27;
13'd2031: Q <= 8'hf2;
13'd2032: Q <= 8'h53;
13'd2033: Q <= 8'hb8;
13'd2034: Q <= 8'h8f;
13'd2035: Q <= 8'ha3;
13'd2036: Q <= 8'h04;
13'd2037: Q <= 8'h23;
13'd2038: Q <= 8'h43;
13'd2039: Q <= 8'h22;
13'd2040: Q <= 8'h17;
13'd2041: Q <= 8'h33;
13'd2042: Q <= 8'h4d;
13'd2043: Q <= 8'h15;
13'd2044: Q <= 8'h50;
13'd2045: Q <= 8'he0;
13'd2046: Q <= 8'h45;
13'd2047: Q <= 8'h00;
13'd2048: Q <= 8'hbf;
13'd2049: Q <= 8'hbe;
13'd2050: Q <= 8'hdf;
13'd2051: Q <= 8'h05;
13'd2052: Q <= 8'h3f;
13'd2053: Q <= 8'h3f;
13'd2054: Q <= 8'h37;
13'd2055: Q <= 8'h08;
13'd2056: Q <= 8'hfa;
13'd2057: Q <= 8'hfd;
13'd2058: Q <= 8'h7f;
13'd2059: Q <= 8'he2;
13'd2060: Q <= 8'hbd;
13'd2061: Q <= 8'hde;
13'd2062: Q <= 8'ha9;
13'd2063: Q <= 8'h0e;
13'd2064: Q <= 8'h98;
13'd2065: Q <= 8'hbc;
13'd2066: Q <= 8'hff;
13'd2067: Q <= 8'hc7;
13'd2068: Q <= 8'h9d;
13'd2069: Q <= 8'h9d;
13'd2070: Q <= 8'h4a;
13'd2071: Q <= 8'h47;
13'd2072: Q <= 8'h9c;
13'd2073: Q <= 8'ha8;
13'd2074: Q <= 8'hfd;
13'd2075: Q <= 8'h24;
13'd2076: Q <= 8'hee;
13'd2077: Q <= 8'haa;
13'd2078: Q <= 8'h9c;
13'd2079: Q <= 8'h80;
13'd2080: Q <= 8'h00;
13'd2081: Q <= 8'h01;
13'd2082: Q <= 8'h00;
13'd2083: Q <= 8'h09;
13'd2084: Q <= 8'h76;
13'd2085: Q <= 8'h1e;
13'd2086: Q <= 8'h8c;
13'd2087: Q <= 8'h84;
13'd2088: Q <= 8'hc9;
13'd2089: Q <= 8'h41;
13'd2090: Q <= 8'h9d;
13'd2091: Q <= 8'h4d;
13'd2092: Q <= 8'h40;
13'd2093: Q <= 8'h08;
13'd2094: Q <= 8'hff;
13'd2095: Q <= 8'hdf;
13'd2096: Q <= 8'ha8;
13'd2097: Q <= 8'h31;
13'd2098: Q <= 8'h1f;
13'd2099: Q <= 8'h3f;
13'd2100: Q <= 8'hba;
13'd2101: Q <= 8'h80;
13'd2102: Q <= 8'h83;
13'd2103: Q <= 8'hc9;
13'd2104: Q <= 8'h91;
13'd2105: Q <= 8'h29;
13'd2106: Q <= 8'h9d;
13'd2107: Q <= 8'hbb;
13'd2108: Q <= 8'h04;
13'd2109: Q <= 8'h00;
13'd2110: Q <= 8'hff;
13'd2111: Q <= 8'h0f;
13'd2112: Q <= 8'ha6;
13'd2113: Q <= 8'h73;
13'd2114: Q <= 8'h04;
13'd2115: Q <= 8'h08;
13'd2116: Q <= 8'ha8;
13'd2117: Q <= 8'h90;
13'd2118: Q <= 8'h00;
13'd2119: Q <= 8'ha0;
13'd2120: Q <= 8'h08;
13'd2121: Q <= 8'h00;
13'd2122: Q <= 8'h00;
13'd2123: Q <= 8'h50;
13'd2124: Q <= 8'h02;
13'd2125: Q <= 8'h00;
13'd2126: Q <= 8'h0c;
13'd2127: Q <= 8'h91;
13'd2128: Q <= 8'hbb;
13'd2129: Q <= 8'h33;
13'd2130: Q <= 8'h08;
13'd2131: Q <= 8'h42;
13'd2132: Q <= 8'h82;
13'd2133: Q <= 8'h00;
13'd2134: Q <= 8'h00;
13'd2135: Q <= 8'ha2;
13'd2136: Q <= 8'h27;
13'd2137: Q <= 8'hb3;
13'd2138: Q <= 8'he1;
13'd2139: Q <= 8'h13;
13'd2140: Q <= 8'h40;
13'd2141: Q <= 8'h10;
13'd2142: Q <= 8'h20;
13'd2143: Q <= 8'h08;
13'd2144: Q <= 8'h00;
13'd2145: Q <= 8'h00;
13'd2146: Q <= 8'h00;
13'd2147: Q <= 8'h00;
13'd2148: Q <= 8'h93;
13'd2149: Q <= 8'h53;
13'd2150: Q <= 8'hcf;
13'd2151: Q <= 8'hc0;
13'd2152: Q <= 8'h4b;
13'd2153: Q <= 8'h1a;
13'd2154: Q <= 8'h07;
13'd2155: Q <= 8'h41;
13'd2156: Q <= 8'h7b;
13'd2157: Q <= 8'h0d;
13'd2158: Q <= 8'h9b;
13'd2159: Q <= 8'h25;
13'd2160: Q <= 8'h0a;
13'd2161: Q <= 8'h02;
13'd2162: Q <= 8'h28;
13'd2163: Q <= 8'h20;
13'd2164: Q <= 8'h00;
13'd2165: Q <= 8'h00;
13'd2166: Q <= 8'h88;
13'd2167: Q <= 8'hd1;
13'd2168: Q <= 8'h27;
13'd2169: Q <= 8'hcc;
13'd2170: Q <= 8'h0a;
13'd2171: Q <= 8'h32;
13'd2172: Q <= 8'h40;
13'd2173: Q <= 8'h01;
13'd2174: Q <= 8'h00;
13'd2175: Q <= 8'h00;
13'd2176: Q <= 8'h10;
13'd2177: Q <= 8'h32;
13'd2178: Q <= 8'h11;
13'd2179: Q <= 8'h10;
13'd2180: Q <= 8'h11;
13'd2181: Q <= 8'h36;
13'd2182: Q <= 8'hfd;
13'd2183: Q <= 8'h10;
13'd2184: Q <= 8'h3d;
13'd2185: Q <= 8'hfd;
13'd2186: Q <= 8'h26;
13'd2187: Q <= 8'h2f;
13'd2188: Q <= 8'hbf;
13'd2189: Q <= 8'h7e;
13'd2190: Q <= 8'h11;
13'd2191: Q <= 8'h01;
13'd2192: Q <= 8'h70;
13'd2193: Q <= 8'hcf;
13'd2194: Q <= 8'hf9;
13'd2195: Q <= 8'hf1;
13'd2196: Q <= 8'hd0;
13'd2197: Q <= 8'h56;
13'd2198: Q <= 8'hf9;
13'd2199: Q <= 8'hb3;
13'd2200: Q <= 8'h00;
13'd2201: Q <= 8'h3b;
13'd2202: Q <= 8'hde;
13'd2203: Q <= 8'haf;
13'd2204: Q <= 8'h18;
13'd2205: Q <= 8'h37;
13'd2206: Q <= 8'h98;
13'd2207: Q <= 8'h39;
13'd2208: Q <= 8'h3f;
13'd2209: Q <= 8'hff;
13'd2210: Q <= 8'hef;
13'd2211: Q <= 8'hfe;
13'd2212: Q <= 8'h82;
13'd2213: Q <= 8'he7;
13'd2214: Q <= 8'h8f;
13'd2215: Q <= 8'h2c;
13'd2216: Q <= 8'h62;
13'd2217: Q <= 8'h80;
13'd2218: Q <= 8'h82;
13'd2219: Q <= 8'hdc;
13'd2220: Q <= 8'h08;
13'd2221: Q <= 8'hf4;
13'd2222: Q <= 8'h18;
13'd2223: Q <= 8'ha8;
13'd2224: Q <= 8'h6f;
13'd2225: Q <= 8'hf0;
13'd2226: Q <= 8'haf;
13'd2227: Q <= 8'hdd;
13'd2228: Q <= 8'ha1;
13'd2229: Q <= 8'he2;
13'd2230: Q <= 8'h5f;
13'd2231: Q <= 8'h64;
13'd2232: Q <= 8'h01;
13'd2233: Q <= 8'h06;
13'd2234: Q <= 8'h03;
13'd2235: Q <= 8'hcc;
13'd2236: Q <= 8'h64;
13'd2237: Q <= 8'hff;
13'd2238: Q <= 8'he4;
13'd2239: Q <= 8'h44;
13'd2240: Q <= 8'h8e;
13'd2241: Q <= 8'h00;
13'd2242: Q <= 8'h10;
13'd2243: Q <= 8'h14;
13'd2244: Q <= 8'h58;
13'd2245: Q <= 8'h10;
13'd2246: Q <= 8'h51;
13'd2247: Q <= 8'h90;
13'd2248: Q <= 8'h45;
13'd2249: Q <= 8'h42;
13'd2250: Q <= 8'h02;
13'd2251: Q <= 8'h31;
13'd2252: Q <= 8'h25;
13'd2253: Q <= 8'h01;
13'd2254: Q <= 8'h35;
13'd2255: Q <= 8'h15;
13'd2256: Q <= 8'h04;
13'd2257: Q <= 8'h28;
13'd2258: Q <= 8'h10;
13'd2259: Q <= 8'h1c;
13'd2260: Q <= 8'h80;
13'd2261: Q <= 8'h00;
13'd2262: Q <= 8'h10;
13'd2263: Q <= 8'h77;
13'd2264: Q <= 8'h5f;
13'd2265: Q <= 8'h8f;
13'd2266: Q <= 8'h02;
13'd2267: Q <= 8'h3f;
13'd2268: Q <= 8'h0c;
13'd2269: Q <= 8'h05;
13'd2270: Q <= 8'h84;
13'd2271: Q <= 8'h3c;
13'd2272: Q <= 8'h21;
13'd2273: Q <= 8'h11;
13'd2274: Q <= 8'hb9;
13'd2275: Q <= 8'h31;
13'd2276: Q <= 8'h00;
13'd2277: Q <= 8'h10;
13'd2278: Q <= 8'h63;
13'd2279: Q <= 8'h23;
13'd2280: Q <= 8'h30;
13'd2281: Q <= 8'h80;
13'd2282: Q <= 8'h33;
13'd2283: Q <= 8'h13;
13'd2284: Q <= 8'h53;
13'd2285: Q <= 8'hd1;
13'd2286: Q <= 8'hbf;
13'd2287: Q <= 8'h15;
13'd2288: Q <= 8'h22;
13'd2289: Q <= 8'h8f;
13'd2290: Q <= 8'haf;
13'd2291: Q <= 8'h38;
13'd2292: Q <= 8'h40;
13'd2293: Q <= 8'h10;
13'd2294: Q <= 8'h02;
13'd2295: Q <= 8'h12;
13'd2296: Q <= 8'h04;
13'd2297: Q <= 8'h90;
13'd2298: Q <= 8'h44;
13'd2299: Q <= 8'h60;
13'd2300: Q <= 8'h64;
13'd2301: Q <= 8'h41;
13'd2302: Q <= 8'hb9;
13'd2303: Q <= 8'h04;
13'd2304: Q <= 8'h20;
13'd2305: Q <= 8'h80;
13'd2306: Q <= 8'h00;
13'd2307: Q <= 8'hb0;
13'd2308: Q <= 8'h00;
13'd2309: Q <= 8'hca;
13'd2310: Q <= 8'h00;
13'd2311: Q <= 8'h80;
13'd2312: Q <= 8'h80;
13'd2313: Q <= 8'h00;
13'd2314: Q <= 8'h00;
13'd2315: Q <= 8'h02;
13'd2316: Q <= 8'h00;
13'd2317: Q <= 8'hbb;
13'd2318: Q <= 8'h00;
13'd2319: Q <= 8'h00;
13'd2320: Q <= 8'h17;
13'd2321: Q <= 8'hbb;
13'd2322: Q <= 8'h00;
13'd2323: Q <= 8'h33;
13'd2324: Q <= 8'h00;
13'd2325: Q <= 8'h00;
13'd2326: Q <= 8'h00;
13'd2327: Q <= 8'h00;
13'd2328: Q <= 8'h20;
13'd2329: Q <= 8'hba;
13'd2330: Q <= 8'h80;
13'd2331: Q <= 8'h89;
13'd2332: Q <= 8'h08;
13'd2333: Q <= 8'haa;
13'd2334: Q <= 8'h00;
13'd2335: Q <= 8'he0;
13'd2336: Q <= 8'hff;
13'd2337: Q <= 8'h0a;
13'd2338: Q <= 8'haf;
13'd2339: Q <= 8'haa;
13'd2340: Q <= 8'h6f;
13'd2341: Q <= 8'h0a;
13'd2342: Q <= 8'hef;
13'd2343: Q <= 8'h0a;
13'd2344: Q <= 8'h02;
13'd2345: Q <= 8'h02;
13'd2346: Q <= 8'h02;
13'd2347: Q <= 8'h20;
13'd2348: Q <= 8'h08;
13'd2349: Q <= 8'h0a;
13'd2350: Q <= 8'h32;
13'd2351: Q <= 8'h08;
13'd2352: Q <= 8'h0e;
13'd2353: Q <= 8'h48;
13'd2354: Q <= 8'hfb;
13'd2355: Q <= 8'ha2;
13'd2356: Q <= 8'h08;
13'd2357: Q <= 8'h10;
13'd2358: Q <= 8'h0b;
13'd2359: Q <= 8'h05;
13'd2360: Q <= 8'h28;
13'd2361: Q <= 8'h00;
13'd2362: Q <= 8'h20;
13'd2363: Q <= 8'h00;
13'd2364: Q <= 8'h00;
13'd2365: Q <= 8'h02;
13'd2366: Q <= 8'h00;
13'd2367: Q <= 8'h00;
13'd2368: Q <= 8'haa;
13'd2369: Q <= 8'hab;
13'd2370: Q <= 8'h10;
13'd2371: Q <= 8'h62;
13'd2372: Q <= 8'he0;
13'd2373: Q <= 8'hc0;
13'd2374: Q <= 8'h80;
13'd2375: Q <= 8'h82;
13'd2376: Q <= 8'h00;
13'd2377: Q <= 8'h00;
13'd2378: Q <= 8'h00;
13'd2379: Q <= 8'h81;
13'd2380: Q <= 8'hc0;
13'd2381: Q <= 8'h80;
13'd2382: Q <= 8'h09;
13'd2383: Q <= 8'ha9;
13'd2384: Q <= 8'hef;
13'd2385: Q <= 8'hba;
13'd2386: Q <= 8'h82;
13'd2387: Q <= 8'h00;
13'd2388: Q <= 8'haa;
13'd2389: Q <= 8'h40;
13'd2390: Q <= 8'h88;
13'd2391: Q <= 8'h02;
13'd2392: Q <= 8'h22;
13'd2393: Q <= 8'h71;
13'd2394: Q <= 8'h03;
13'd2395: Q <= 8'h02;
13'd2396: Q <= 8'h80;
13'd2397: Q <= 8'h80;
13'd2398: Q <= 8'h40;
13'd2399: Q <= 8'h01;
13'd2400: Q <= 8'h5d;
13'd2401: Q <= 8'h31;
13'd2402: Q <= 8'h80;
13'd2403: Q <= 8'h24;
13'd2404: Q <= 8'h59;
13'd2405: Q <= 8'h00;
13'd2406: Q <= 8'h26;
13'd2407: Q <= 8'h1e;
13'd2408: Q <= 8'hfb;
13'd2409: Q <= 8'h19;
13'd2410: Q <= 8'h94;
13'd2411: Q <= 8'h15;
13'd2412: Q <= 8'h11;
13'd2413: Q <= 8'h01;
13'd2414: Q <= 8'h00;
13'd2415: Q <= 8'h1b;
13'd2416: Q <= 8'hba;
13'd2417: Q <= 8'hc9;
13'd2418: Q <= 8'h8e;
13'd2419: Q <= 8'hef;
13'd2420: Q <= 8'he8;
13'd2421: Q <= 8'h89;
13'd2422: Q <= 8'h88;
13'd2423: Q <= 8'h8d;
13'd2424: Q <= 8'hf0;
13'd2425: Q <= 8'h44;
13'd2426: Q <= 8'hc0;
13'd2427: Q <= 8'h00;
13'd2428: Q <= 8'h00;
13'd2429: Q <= 8'h10;
13'd2430: Q <= 8'h00;
13'd2431: Q <= 8'h08;
13'd2432: Q <= 8'h20;
13'd2433: Q <= 8'h12;
13'd2434: Q <= 8'h04;
13'd2435: Q <= 8'h30;
13'd2436: Q <= 8'ha0;
13'd2437: Q <= 8'h00;
13'd2438: Q <= 8'h00;
13'd2439: Q <= 8'h00;
13'd2440: Q <= 8'h06;
13'd2441: Q <= 8'h01;
13'd2442: Q <= 8'h08;
13'd2443: Q <= 8'h21;
13'd2444: Q <= 8'hbf;
13'd2445: Q <= 8'h15;
13'd2446: Q <= 8'h9f;
13'd2447: Q <= 8'h1f;
13'd2448: Q <= 8'hb0;
13'd2449: Q <= 8'h08;
13'd2450: Q <= 8'h00;
13'd2451: Q <= 8'h01;
13'd2452: Q <= 8'h88;
13'd2453: Q <= 8'h00;
13'd2454: Q <= 8'hc0;
13'd2455: Q <= 8'h88;
13'd2456: Q <= 8'hb2;
13'd2457: Q <= 8'hc2;
13'd2458: Q <= 8'h00;
13'd2459: Q <= 8'h02;
13'd2460: Q <= 8'h88;
13'd2461: Q <= 8'h08;
13'd2462: Q <= 8'h00;
13'd2463: Q <= 8'h09;
13'd2464: Q <= 8'hcf;
13'd2465: Q <= 8'he7;
13'd2466: Q <= 8'hff;
13'd2467: Q <= 8'hff;
13'd2468: Q <= 8'h0c;
13'd2469: Q <= 8'he4;
13'd2470: Q <= 8'h0f;
13'd2471: Q <= 8'he6;
13'd2472: Q <= 8'h02;
13'd2473: Q <= 8'h80;
13'd2474: Q <= 8'h88;
13'd2475: Q <= 8'ha8;
13'd2476: Q <= 8'h4e;
13'd2477: Q <= 8'hf7;
13'd2478: Q <= 8'h01;
13'd2479: Q <= 8'h86;
13'd2480: Q <= 8'hce;
13'd2481: Q <= 8'haa;
13'd2482: Q <= 8'hdf;
13'd2483: Q <= 8'h5f;
13'd2484: Q <= 8'h10;
13'd2485: Q <= 8'h91;
13'd2486: Q <= 8'h48;
13'd2487: Q <= 8'h00;
13'd2488: Q <= 8'h00;
13'd2489: Q <= 8'hc0;
13'd2490: Q <= 8'h8f;
13'd2491: Q <= 8'h40;
13'd2492: Q <= 8'h04;
13'd2493: Q <= 8'hf4;
13'd2494: Q <= 8'h40;
13'd2495: Q <= 8'h04;
13'd2496: Q <= 8'h7e;
13'd2497: Q <= 8'h20;
13'd2498: Q <= 8'h7c;
13'd2499: Q <= 8'h02;
13'd2500: Q <= 8'h89;
13'd2501: Q <= 8'h10;
13'd2502: Q <= 8'h32;
13'd2503: Q <= 8'h00;
13'd2504: Q <= 8'h70;
13'd2505: Q <= 8'h00;
13'd2506: Q <= 8'h88;
13'd2507: Q <= 8'h91;
13'd2508: Q <= 8'hba;
13'd2509: Q <= 8'h90;
13'd2510: Q <= 8'h13;
13'd2511: Q <= 8'h19;
13'd2512: Q <= 8'h40;
13'd2513: Q <= 8'h80;
13'd2514: Q <= 8'hca;
13'd2515: Q <= 8'h18;
13'd2516: Q <= 8'hb7;
13'd2517: Q <= 8'h10;
13'd2518: Q <= 8'h1b;
13'd2519: Q <= 8'h10;
13'd2520: Q <= 8'hf8;
13'd2521: Q <= 8'h08;
13'd2522: Q <= 8'hde;
13'd2523: Q <= 8'h40;
13'd2524: Q <= 8'hff;
13'd2525: Q <= 8'h3f;
13'd2526: Q <= 8'h31;
13'd2527: Q <= 8'h31;
13'd2528: Q <= 8'h0b;
13'd2529: Q <= 8'h3f;
13'd2530: Q <= 8'hff;
13'd2531: Q <= 8'h06;
13'd2532: Q <= 8'h03;
13'd2533: Q <= 8'hf9;
13'd2534: Q <= 8'h83;
13'd2535: Q <= 8'h02;
13'd2536: Q <= 8'h42;
13'd2537: Q <= 8'h01;
13'd2538: Q <= 8'h00;
13'd2539: Q <= 8'h84;
13'd2540: Q <= 8'h24;
13'd2541: Q <= 8'he1;
13'd2542: Q <= 8'h02;
13'd2543: Q <= 8'h00;
13'd2544: Q <= 8'h64;
13'd2545: Q <= 8'h63;
13'd2546: Q <= 8'h4e;
13'd2547: Q <= 8'h20;
13'd2548: Q <= 8'hc3;
13'd2549: Q <= 8'hd2;
13'd2550: Q <= 8'h44;
13'd2551: Q <= 8'h15;
13'd2552: Q <= 8'h60;
13'd2553: Q <= 8'h40;
13'd2554: Q <= 8'h09;
13'd2555: Q <= 8'h41;
13'd2556: Q <= 8'h20;
13'd2557: Q <= 8'hd7;
13'd2558: Q <= 8'h00;
13'd2559: Q <= 8'h40;
13'd2560: Q <= 8'h60;
13'd2561: Q <= 8'h17;
13'd2562: Q <= 8'h80;
13'd2563: Q <= 8'h10;
13'd2564: Q <= 8'h97;
13'd2565: Q <= 8'h7c;
13'd2566: Q <= 8'hd2;
13'd2567: Q <= 8'had;
13'd2568: Q <= 8'h3e;
13'd2569: Q <= 8'h12;
13'd2570: Q <= 8'h00;
13'd2571: Q <= 8'h50;
13'd2572: Q <= 8'hdd;
13'd2573: Q <= 8'hf1;
13'd2574: Q <= 8'hdc;
13'd2575: Q <= 8'hd2;
13'd2576: Q <= 8'hc0;
13'd2577: Q <= 8'h04;
13'd2578: Q <= 8'h00;
13'd2579: Q <= 8'hc0;
13'd2580: Q <= 8'hc8;
13'd2581: Q <= 8'h04;
13'd2582: Q <= 8'hd2;
13'd2583: Q <= 8'h10;
13'd2584: Q <= 8'h8c;
13'd2585: Q <= 8'h04;
13'd2586: Q <= 8'hc8;
13'd2587: Q <= 8'h18;
13'd2588: Q <= 8'hdc;
13'd2589: Q <= 8'h51;
13'd2590: Q <= 8'hd0;
13'd2591: Q <= 8'hf5;
13'd2592: Q <= 8'h30;
13'd2593: Q <= 8'h27;
13'd2594: Q <= 8'h73;
13'd2595: Q <= 8'h2f;
13'd2596: Q <= 8'h80;
13'd2597: Q <= 8'h60;
13'd2598: Q <= 8'h57;
13'd2599: Q <= 8'h07;
13'd2600: Q <= 8'h10;
13'd2601: Q <= 8'h00;
13'd2602: Q <= 8'h04;
13'd2603: Q <= 8'h82;
13'd2604: Q <= 8'h34;
13'd2605: Q <= 8'h40;
13'd2606: Q <= 8'hf7;
13'd2607: Q <= 8'h0c;
13'd2608: Q <= 8'h01;
13'd2609: Q <= 8'h13;
13'd2610: Q <= 8'h02;
13'd2611: Q <= 8'h42;
13'd2612: Q <= 8'h00;
13'd2613: Q <= 8'h40;
13'd2614: Q <= 8'h00;
13'd2615: Q <= 8'h00;
13'd2616: Q <= 8'h00;
13'd2617: Q <= 8'h13;
13'd2618: Q <= 8'h10;
13'd2619: Q <= 8'h30;
13'd2620: Q <= 8'h22;
13'd2621: Q <= 8'h11;
13'd2622: Q <= 8'h51;
13'd2623: Q <= 8'h17;
13'd2624: Q <= 8'hdd;
13'd2625: Q <= 8'h15;
13'd2626: Q <= 8'h10;
13'd2627: Q <= 8'h35;
13'd2628: Q <= 8'h04;
13'd2629: Q <= 8'h18;
13'd2630: Q <= 8'h13;
13'd2631: Q <= 8'hff;
13'd2632: Q <= 8'hf5;
13'd2633: Q <= 8'h90;
13'd2634: Q <= 8'h11;
13'd2635: Q <= 8'h1d;
13'd2636: Q <= 8'h31;
13'd2637: Q <= 8'h10;
13'd2638: Q <= 8'h31;
13'd2639: Q <= 8'hfd;
13'd2640: Q <= 8'h9a;
13'd2641: Q <= 8'h88;
13'd2642: Q <= 8'h42;
13'd2643: Q <= 8'h48;
13'd2644: Q <= 8'h00;
13'd2645: Q <= 8'h08;
13'd2646: Q <= 8'h00;
13'd2647: Q <= 8'h4d;
13'd2648: Q <= 8'h91;
13'd2649: Q <= 8'h09;
13'd2650: Q <= 8'h10;
13'd2651: Q <= 8'h04;
13'd2652: Q <= 8'h20;
13'd2653: Q <= 8'h09;
13'd2654: Q <= 8'h01;
13'd2655: Q <= 8'h1c;
13'd2656: Q <= 8'h0c;
13'd2657: Q <= 8'hf8;
13'd2658: Q <= 8'h21;
13'd2659: Q <= 8'h51;
13'd2660: Q <= 8'h08;
13'd2661: Q <= 8'h51;
13'd2662: Q <= 8'h21;
13'd2663: Q <= 8'h71;
13'd2664: Q <= 8'h8a;
13'd2665: Q <= 8'h10;
13'd2666: Q <= 8'h01;
13'd2667: Q <= 8'h41;
13'd2668: Q <= 8'h16;
13'd2669: Q <= 8'h03;
13'd2670: Q <= 8'h03;
13'd2671: Q <= 8'h11;
13'd2672: Q <= 8'h08;
13'd2673: Q <= 8'h30;
13'd2674: Q <= 8'h04;
13'd2675: Q <= 8'h40;
13'd2676: Q <= 8'h00;
13'd2677: Q <= 8'h28;
13'd2678: Q <= 8'h18;
13'd2679: Q <= 8'h32;
13'd2680: Q <= 8'h10;
13'd2681: Q <= 8'h00;
13'd2682: Q <= 8'h04;
13'd2683: Q <= 8'h80;
13'd2684: Q <= 8'h00;
13'd2685: Q <= 8'h00;
13'd2686: Q <= 8'h04;
13'd2687: Q <= 8'h00;
13'd2688: Q <= 8'hfb;
13'd2689: Q <= 8'h0e;
13'd2690: Q <= 8'hfe;
13'd2691: Q <= 8'haa;
13'd2692: Q <= 8'h50;
13'd2693: Q <= 8'h00;
13'd2694: Q <= 8'hca;
13'd2695: Q <= 8'h8e;
13'd2696: Q <= 8'hec;
13'd2697: Q <= 8'h81;
13'd2698: Q <= 8'h48;
13'd2699: Q <= 8'h80;
13'd2700: Q <= 8'h90;
13'd2701: Q <= 8'h04;
13'd2702: Q <= 8'h80;
13'd2703: Q <= 8'h08;
13'd2704: Q <= 8'h03;
13'd2705: Q <= 8'h03;
13'd2706: Q <= 8'h4b;
13'd2707: Q <= 8'h1e;
13'd2708: Q <= 8'h00;
13'd2709: Q <= 8'h08;
13'd2710: Q <= 8'h49;
13'd2711: Q <= 8'h01;
13'd2712: Q <= 8'h40;
13'd2713: Q <= 8'h42;
13'd2714: Q <= 8'h80;
13'd2715: Q <= 8'h02;
13'd2716: Q <= 8'h40;
13'd2717: Q <= 8'h00;
13'd2718: Q <= 8'h00;
13'd2719: Q <= 8'h00;
13'd2720: Q <= 8'h6c;
13'd2721: Q <= 8'h2c;
13'd2722: Q <= 8'h00;
13'd2723: Q <= 8'h0c;
13'd2724: Q <= 8'hdd;
13'd2725: Q <= 8'h1c;
13'd2726: Q <= 8'h5f;
13'd2727: Q <= 8'hff;
13'd2728: Q <= 8'haf;
13'd2729: Q <= 8'hac;
13'd2730: Q <= 8'h18;
13'd2731: Q <= 8'h0e;
13'd2732: Q <= 8'h8c;
13'd2733: Q <= 8'h0a;
13'd2734: Q <= 8'h7a;
13'd2735: Q <= 8'h2c;
13'd2736: Q <= 8'h3e;
13'd2737: Q <= 8'h84;
13'd2738: Q <= 8'h4e;
13'd2739: Q <= 8'h8a;
13'd2740: Q <= 8'h3e;
13'd2741: Q <= 8'h00;
13'd2742: Q <= 8'he8;
13'd2743: Q <= 8'h00;
13'd2744: Q <= 8'h4e;
13'd2745: Q <= 8'hce;
13'd2746: Q <= 8'h0c;
13'd2747: Q <= 8'hc9;
13'd2748: Q <= 8'h44;
13'd2749: Q <= 8'h0f;
13'd2750: Q <= 8'h54;
13'd2751: Q <= 8'h0b;
13'd2752: Q <= 8'h2b;
13'd2753: Q <= 8'h63;
13'd2754: Q <= 8'h77;
13'd2755: Q <= 8'h23;
13'd2756: Q <= 8'h07;
13'd2757: Q <= 8'he6;
13'd2758: Q <= 8'h1f;
13'd2759: Q <= 8'h27;
13'd2760: Q <= 8'h12;
13'd2761: Q <= 8'h43;
13'd2762: Q <= 8'h03;
13'd2763: Q <= 8'h10;
13'd2764: Q <= 8'h8a;
13'd2765: Q <= 8'h41;
13'd2766: Q <= 8'h10;
13'd2767: Q <= 8'h22;
13'd2768: Q <= 8'h47;
13'd2769: Q <= 8'h07;
13'd2770: Q <= 8'h43;
13'd2771: Q <= 8'h1a;
13'd2772: Q <= 8'h0a;
13'd2773: Q <= 8'h08;
13'd2774: Q <= 8'h02;
13'd2775: Q <= 8'h00;
13'd2776: Q <= 8'h47;
13'd2777: Q <= 8'h05;
13'd2778: Q <= 8'h63;
13'd2779: Q <= 8'h15;
13'd2780: Q <= 8'h45;
13'd2781: Q <= 8'hf7;
13'd2782: Q <= 8'h73;
13'd2783: Q <= 8'h77;
13'd2784: Q <= 8'h0b;
13'd2785: Q <= 8'h2f;
13'd2786: Q <= 8'hdf;
13'd2787: Q <= 8'hc7;
13'd2788: Q <= 8'h81;
13'd2789: Q <= 8'hf0;
13'd2790: Q <= 8'h08;
13'd2791: Q <= 8'h42;
13'd2792: Q <= 8'h8a;
13'd2793: Q <= 8'h40;
13'd2794: Q <= 8'h8f;
13'd2795: Q <= 8'hb0;
13'd2796: Q <= 8'h06;
13'd2797: Q <= 8'he2;
13'd2798: Q <= 8'h08;
13'd2799: Q <= 8'h04;
13'd2800: Q <= 8'h4c;
13'd2801: Q <= 8'h07;
13'd2802: Q <= 8'h17;
13'd2803: Q <= 8'h51;
13'd2804: Q <= 8'h4d;
13'd2805: Q <= 8'h05;
13'd2806: Q <= 8'hc8;
13'd2807: Q <= 8'h5c;
13'd2808: Q <= 8'h41;
13'd2809: Q <= 8'h42;
13'd2810: Q <= 8'h4e;
13'd2811: Q <= 8'h24;
13'd2812: Q <= 8'h4a;
13'd2813: Q <= 8'hf6;
13'd2814: Q <= 8'h46;
13'd2815: Q <= 8'hd4;
13'd2816: Q <= 8'h40;
13'd2817: Q <= 8'h27;
13'd2818: Q <= 8'h05;
13'd2819: Q <= 8'h01;
13'd2820: Q <= 8'h21;
13'd2821: Q <= 8'h0c;
13'd2822: Q <= 8'h4f;
13'd2823: Q <= 8'h0e;
13'd2824: Q <= 8'h79;
13'd2825: Q <= 8'h0f;
13'd2826: Q <= 8'h71;
13'd2827: Q <= 8'ha3;
13'd2828: Q <= 8'h33;
13'd2829: Q <= 8'h0e;
13'd2830: Q <= 8'hef;
13'd2831: Q <= 8'h04;
13'd2832: Q <= 8'h73;
13'd2833: Q <= 8'h33;
13'd2834: Q <= 8'h93;
13'd2835: Q <= 8'h37;
13'd2836: Q <= 8'h78;
13'd2837: Q <= 8'hcf;
13'd2838: Q <= 8'hfe;
13'd2839: Q <= 8'h4d;
13'd2840: Q <= 8'h55;
13'd2841: Q <= 8'h5f;
13'd2842: Q <= 8'hbf;
13'd2843: Q <= 8'h1f;
13'd2844: Q <= 8'h34;
13'd2845: Q <= 8'h44;
13'd2846: Q <= 8'he7;
13'd2847: Q <= 8'h05;
13'd2848: Q <= 8'hd5;
13'd2849: Q <= 8'h54;
13'd2850: Q <= 8'h18;
13'd2851: Q <= 8'h27;
13'd2852: Q <= 8'h74;
13'd2853: Q <= 8'hbb;
13'd2854: Q <= 8'h39;
13'd2855: Q <= 8'hac;
13'd2856: Q <= 8'h2b;
13'd2857: Q <= 8'h22;
13'd2858: Q <= 8'hfb;
13'd2859: Q <= 8'h37;
13'd2860: Q <= 8'h33;
13'd2861: Q <= 8'h43;
13'd2862: Q <= 8'ha6;
13'd2863: Q <= 8'h8f;
13'd2864: Q <= 8'hd5;
13'd2865: Q <= 8'hfc;
13'd2866: Q <= 8'hbb;
13'd2867: Q <= 8'h1d;
13'd2868: Q <= 8'hf2;
13'd2869: Q <= 8'hf7;
13'd2870: Q <= 8'ha7;
13'd2871: Q <= 8'hde;
13'd2872: Q <= 8'h54;
13'd2873: Q <= 8'h7b;
13'd2874: Q <= 8'hf3;
13'd2875: Q <= 8'h72;
13'd2876: Q <= 8'h40;
13'd2877: Q <= 8'h0c;
13'd2878: Q <= 8'h10;
13'd2879: Q <= 8'h11;
13'd2880: Q <= 8'h50;
13'd2881: Q <= 8'h7a;
13'd2882: Q <= 8'h04;
13'd2883: Q <= 8'h14;
13'd2884: Q <= 8'h50;
13'd2885: Q <= 8'h51;
13'd2886: Q <= 8'h18;
13'd2887: Q <= 8'h91;
13'd2888: Q <= 8'h59;
13'd2889: Q <= 8'h00;
13'd2890: Q <= 8'h00;
13'd2891: Q <= 8'h00;
13'd2892: Q <= 8'hf1;
13'd2893: Q <= 8'h71;
13'd2894: Q <= 8'h00;
13'd2895: Q <= 8'h74;
13'd2896: Q <= 8'h88;
13'd2897: Q <= 8'h99;
13'd2898: Q <= 8'h80;
13'd2899: Q <= 8'hc8;
13'd2900: Q <= 8'hc4;
13'd2901: Q <= 8'hb0;
13'd2902: Q <= 8'h00;
13'd2903: Q <= 8'hf1;
13'd2904: Q <= 8'h02;
13'd2905: Q <= 8'h00;
13'd2906: Q <= 8'h00;
13'd2907: Q <= 8'h88;
13'd2908: Q <= 8'hc4;
13'd2909: Q <= 8'h30;
13'd2910: Q <= 8'h02;
13'd2911: Q <= 8'h28;
13'd2912: Q <= 8'h2f;
13'd2913: Q <= 8'haf;
13'd2914: Q <= 8'hbf;
13'd2915: Q <= 8'hfd;
13'd2916: Q <= 8'h87;
13'd2917: Q <= 8'h3e;
13'd2918: Q <= 8'h36;
13'd2919: Q <= 8'h08;
13'd2920: Q <= 8'h32;
13'd2921: Q <= 8'ha6;
13'd2922: Q <= 8'haa;
13'd2923: Q <= 8'he9;
13'd2924: Q <= 8'h96;
13'd2925: Q <= 8'hbc;
13'd2926: Q <= 8'ha1;
13'd2927: Q <= 8'h88;
13'd2928: Q <= 8'h41;
13'd2929: Q <= 8'h66;
13'd2930: Q <= 8'hf5;
13'd2931: Q <= 8'h1f;
13'd2932: Q <= 8'h77;
13'd2933: Q <= 8'hd8;
13'd2934: Q <= 8'h04;
13'd2935: Q <= 8'h62;
13'd2936: Q <= 8'h04;
13'd2937: Q <= 8'h05;
13'd2938: Q <= 8'he6;
13'd2939: Q <= 8'hcf;
13'd2940: Q <= 8'h75;
13'd2941: Q <= 8'hfb;
13'd2942: Q <= 8'h46;
13'd2943: Q <= 8'hc0;
13'd2944: Q <= 8'h80;
13'd2945: Q <= 8'h15;
13'd2946: Q <= 8'h00;
13'd2947: Q <= 8'h00;
13'd2948: Q <= 8'h00;
13'd2949: Q <= 8'h51;
13'd2950: Q <= 8'h00;
13'd2951: Q <= 8'h80;
13'd2952: Q <= 8'h45;
13'd2953: Q <= 8'h5d;
13'd2954: Q <= 8'h40;
13'd2955: Q <= 8'h80;
13'd2956: Q <= 8'h5d;
13'd2957: Q <= 8'hd5;
13'd2958: Q <= 8'h44;
13'd2959: Q <= 8'h00;
13'd2960: Q <= 8'h41;
13'd2961: Q <= 8'h40;
13'd2962: Q <= 8'h00;
13'd2963: Q <= 8'h00;
13'd2964: Q <= 8'h00;
13'd2965: Q <= 8'h01;
13'd2966: Q <= 8'h00;
13'd2967: Q <= 8'h00;
13'd2968: Q <= 8'h57;
13'd2969: Q <= 8'h55;
13'd2970: Q <= 8'h00;
13'd2971: Q <= 8'h0c;
13'd2972: Q <= 8'h55;
13'd2973: Q <= 8'h75;
13'd2974: Q <= 8'h40;
13'd2975: Q <= 8'h04;
13'd2976: Q <= 8'h1b;
13'd2977: Q <= 8'h0c;
13'd2978: Q <= 8'h28;
13'd2979: Q <= 8'h08;
13'd2980: Q <= 8'hb4;
13'd2981: Q <= 8'h2e;
13'd2982: Q <= 8'hc3;
13'd2983: Q <= 8'h1d;
13'd2984: Q <= 8'hdb;
13'd2985: Q <= 8'hb5;
13'd2986: Q <= 8'he1;
13'd2987: Q <= 8'h87;
13'd2988: Q <= 8'h35;
13'd2989: Q <= 8'h26;
13'd2990: Q <= 8'h31;
13'd2991: Q <= 8'h05;
13'd2992: Q <= 8'hcf;
13'd2993: Q <= 8'h0a;
13'd2994: Q <= 8'h3f;
13'd2995: Q <= 8'h26;
13'd2996: Q <= 8'h5e;
13'd2997: Q <= 8'hee;
13'd2998: Q <= 8'hff;
13'd2999: Q <= 8'h2e;
13'd3000: Q <= 8'hd7;
13'd3001: Q <= 8'h06;
13'd3002: Q <= 8'h6b;
13'd3003: Q <= 8'h44;
13'd3004: Q <= 8'h12;
13'd3005: Q <= 8'h4c;
13'd3006: Q <= 8'h0a;
13'd3007: Q <= 8'h08;
13'd3008: Q <= 8'hef;
13'd3009: Q <= 8'h00;
13'd3010: Q <= 8'hc0;
13'd3011: Q <= 8'h08;
13'd3012: Q <= 8'haa;
13'd3013: Q <= 8'h44;
13'd3014: Q <= 8'h1e;
13'd3015: Q <= 8'h6a;
13'd3016: Q <= 8'h0e;
13'd3017: Q <= 8'h1a;
13'd3018: Q <= 8'h2a;
13'd3019: Q <= 8'h82;
13'd3020: Q <= 8'heb;
13'd3021: Q <= 8'h08;
13'd3022: Q <= 8'h66;
13'd3023: Q <= 8'h08;
13'd3024: Q <= 8'h4e;
13'd3025: Q <= 8'h01;
13'd3026: Q <= 8'h00;
13'd3027: Q <= 8'h01;
13'd3028: Q <= 8'h1c;
13'd3029: Q <= 8'h02;
13'd3030: Q <= 8'h08;
13'd3031: Q <= 8'h74;
13'd3032: Q <= 8'h6a;
13'd3033: Q <= 8'h0a;
13'd3034: Q <= 8'h23;
13'd3035: Q <= 8'h62;
13'd3036: Q <= 8'h2a;
13'd3037: Q <= 8'h23;
13'd3038: Q <= 8'h04;
13'd3039: Q <= 8'h32;
13'd3040: Q <= 8'h11;
13'd3041: Q <= 8'h23;
13'd3042: Q <= 8'h98;
13'd3043: Q <= 8'h31;
13'd3044: Q <= 8'h12;
13'd3045: Q <= 8'h00;
13'd3046: Q <= 8'h83;
13'd3047: Q <= 8'h3a;
13'd3048: Q <= 8'h88;
13'd3049: Q <= 8'h01;
13'd3050: Q <= 8'h00;
13'd3051: Q <= 8'h12;
13'd3052: Q <= 8'h80;
13'd3053: Q <= 8'h00;
13'd3054: Q <= 8'h80;
13'd3055: Q <= 8'h22;
13'd3056: Q <= 8'h17;
13'd3057: Q <= 8'h0f;
13'd3058: Q <= 8'h92;
13'd3059: Q <= 8'h37;
13'd3060: Q <= 8'h02;
13'd3061: Q <= 8'h02;
13'd3062: Q <= 8'h0e;
13'd3063: Q <= 8'h77;
13'd3064: Q <= 8'h00;
13'd3065: Q <= 8'h03;
13'd3066: Q <= 8'h00;
13'd3067: Q <= 8'h02;
13'd3068: Q <= 8'h00;
13'd3069: Q <= 8'h00;
13'd3070: Q <= 8'h20;
13'd3071: Q <= 8'h04;
13'd3072: Q <= 8'h00;
13'd3073: Q <= 8'h0d;
13'd3074: Q <= 8'h10;
13'd3075: Q <= 8'h07;
13'd3076: Q <= 8'h08;
13'd3077: Q <= 8'h49;
13'd3078: Q <= 8'h10;
13'd3079: Q <= 8'h48;
13'd3080: Q <= 8'h21;
13'd3081: Q <= 8'h0d;
13'd3082: Q <= 8'h4d;
13'd3083: Q <= 8'hbd;
13'd3084: Q <= 8'h88;
13'd3085: Q <= 8'h01;
13'd3086: Q <= 8'h88;
13'd3087: Q <= 8'h4f;
13'd3088: Q <= 8'hfd;
13'd3089: Q <= 8'hbf;
13'd3090: Q <= 8'ha9;
13'd3091: Q <= 8'hbd;
13'd3092: Q <= 8'h90;
13'd3093: Q <= 8'hbb;
13'd3094: Q <= 8'hb8;
13'd3095: Q <= 8'h11;
13'd3096: Q <= 8'h84;
13'd3097: Q <= 8'hd9;
13'd3098: Q <= 8'hcf;
13'd3099: Q <= 8'had;
13'd3100: Q <= 8'h88;
13'd3101: Q <= 8'h21;
13'd3102: Q <= 8'h50;
13'd3103: Q <= 8'h08;
13'd3104: Q <= 8'h23;
13'd3105: Q <= 8'h67;
13'd3106: Q <= 8'h2f;
13'd3107: Q <= 8'h66;
13'd3108: Q <= 8'h27;
13'd3109: Q <= 8'hea;
13'd3110: Q <= 8'h23;
13'd3111: Q <= 8'h00;
13'd3112: Q <= 8'hee;
13'd3113: Q <= 8'h6e;
13'd3114: Q <= 8'hae;
13'd3115: Q <= 8'h06;
13'd3116: Q <= 8'h23;
13'd3117: Q <= 8'h6e;
13'd3118: Q <= 8'hc2;
13'd3119: Q <= 8'h20;
13'd3120: Q <= 8'h47;
13'd3121: Q <= 8'h6b;
13'd3122: Q <= 8'h67;
13'd3123: Q <= 8'h5d;
13'd3124: Q <= 8'hbf;
13'd3125: Q <= 8'hff;
13'd3126: Q <= 8'h6e;
13'd3127: Q <= 8'h66;
13'd3128: Q <= 8'h03;
13'd3129: Q <= 8'h50;
13'd3130: Q <= 8'h67;
13'd3131: Q <= 8'h14;
13'd3132: Q <= 8'h42;
13'd3133: Q <= 8'hc6;
13'd3134: Q <= 8'h12;
13'd3135: Q <= 8'h40;
13'd3136: Q <= 8'h75;
13'd3137: Q <= 8'h59;
13'd3138: Q <= 8'h14;
13'd3139: Q <= 8'h05;
13'd3140: Q <= 8'hd5;
13'd3141: Q <= 8'h75;
13'd3142: Q <= 8'h1d;
13'd3143: Q <= 8'hed;
13'd3144: Q <= 8'hfe;
13'd3145: Q <= 8'h81;
13'd3146: Q <= 8'h00;
13'd3147: Q <= 8'h00;
13'd3148: Q <= 8'hcf;
13'd3149: Q <= 8'h75;
13'd3150: Q <= 8'h74;
13'd3151: Q <= 8'h8e;
13'd3152: Q <= 8'h8c;
13'd3153: Q <= 8'h10;
13'd3154: Q <= 8'hcd;
13'd3155: Q <= 8'h81;
13'd3156: Q <= 8'h88;
13'd3157: Q <= 8'h0b;
13'd3158: Q <= 8'h8d;
13'd3159: Q <= 8'h0f;
13'd3160: Q <= 8'hfe;
13'd3161: Q <= 8'hc0;
13'd3162: Q <= 8'h0a;
13'd3163: Q <= 8'h25;
13'd3164: Q <= 8'h19;
13'd3165: Q <= 8'h0c;
13'd3166: Q <= 8'h48;
13'd3167: Q <= 8'h05;
13'd3168: Q <= 8'h58;
13'd3169: Q <= 8'h10;
13'd3170: Q <= 8'h90;
13'd3171: Q <= 8'h11;
13'd3172: Q <= 8'h00;
13'd3173: Q <= 8'h90;
13'd3174: Q <= 8'h13;
13'd3175: Q <= 8'h15;
13'd3176: Q <= 8'h05;
13'd3177: Q <= 8'h1c;
13'd3178: Q <= 8'hd2;
13'd3179: Q <= 8'h61;
13'd3180: Q <= 8'h10;
13'd3181: Q <= 8'h01;
13'd3182: Q <= 8'h00;
13'd3183: Q <= 8'h03;
13'd3184: Q <= 8'h24;
13'd3185: Q <= 8'h03;
13'd3186: Q <= 8'h08;
13'd3187: Q <= 8'h7c;
13'd3188: Q <= 8'h00;
13'd3189: Q <= 8'h00;
13'd3190: Q <= 8'hb8;
13'd3191: Q <= 8'hbb;
13'd3192: Q <= 8'h28;
13'd3193: Q <= 8'h08;
13'd3194: Q <= 8'h88;
13'd3195: Q <= 8'h08;
13'd3196: Q <= 8'h04;
13'd3197: Q <= 8'h02;
13'd3198: Q <= 8'h10;
13'd3199: Q <= 8'h09;
13'd3200: Q <= 8'h25;
13'd3201: Q <= 8'hbe;
13'd3202: Q <= 8'h7f;
13'd3203: Q <= 8'h8f;
13'd3204: Q <= 8'h2f;
13'd3205: Q <= 8'h6f;
13'd3206: Q <= 8'h0f;
13'd3207: Q <= 8'h26;
13'd3208: Q <= 8'hf2;
13'd3209: Q <= 8'ha6;
13'd3210: Q <= 8'hef;
13'd3211: Q <= 8'h6f;
13'd3212: Q <= 8'h4b;
13'd3213: Q <= 8'hb2;
13'd3214: Q <= 8'h0b;
13'd3215: Q <= 8'h02;
13'd3216: Q <= 8'h4e;
13'd3217: Q <= 8'h33;
13'd3218: Q <= 8'hd7;
13'd3219: Q <= 8'h3f;
13'd3220: Q <= 8'h87;
13'd3221: Q <= 8'h54;
13'd3222: Q <= 8'h6b;
13'd3223: Q <= 8'h27;
13'd3224: Q <= 8'h24;
13'd3225: Q <= 8'h09;
13'd3226: Q <= 8'hc5;
13'd3227: Q <= 8'h22;
13'd3228: Q <= 8'h9e;
13'd3229: Q <= 8'hc6;
13'd3230: Q <= 8'hce;
13'd3231: Q <= 8'hc0;
13'd3232: Q <= 8'hbf;
13'd3233: Q <= 8'h33;
13'd3234: Q <= 8'h40;
13'd3235: Q <= 8'h3b;
13'd3236: Q <= 8'h09;
13'd3237: Q <= 8'h10;
13'd3238: Q <= 8'h1b;
13'd3239: Q <= 8'hbf;
13'd3240: Q <= 8'h7b;
13'd3241: Q <= 8'h11;
13'd3242: Q <= 8'h01;
13'd3243: Q <= 8'h13;
13'd3244: Q <= 8'ha0;
13'd3245: Q <= 8'h00;
13'd3246: Q <= 8'h11;
13'd3247: Q <= 8'h13;
13'd3248: Q <= 8'h2a;
13'd3249: Q <= 8'h2b;
13'd3250: Q <= 8'h48;
13'd3251: Q <= 8'hbe;
13'd3252: Q <= 8'h48;
13'd3253: Q <= 8'h08;
13'd3254: Q <= 8'h88;
13'd3255: Q <= 8'hba;
13'd3256: Q <= 8'h4d;
13'd3257: Q <= 8'haf;
13'd3258: Q <= 8'h40;
13'd3259: Q <= 8'h07;
13'd3260: Q <= 8'h40;
13'd3261: Q <= 8'h08;
13'd3262: Q <= 8'h08;
13'd3263: Q <= 8'h08;
13'd3264: Q <= 8'h50;
13'd3265: Q <= 8'h50;
13'd3266: Q <= 8'h00;
13'd3267: Q <= 8'h11;
13'd3268: Q <= 8'h0a;
13'd3269: Q <= 8'h61;
13'd3270: Q <= 8'h20;
13'd3271: Q <= 8'h20;
13'd3272: Q <= 8'h20;
13'd3273: Q <= 8'h10;
13'd3274: Q <= 8'h00;
13'd3275: Q <= 8'h94;
13'd3276: Q <= 8'h54;
13'd3277: Q <= 8'h10;
13'd3278: Q <= 8'h02;
13'd3279: Q <= 8'h16;
13'd3280: Q <= 8'h10;
13'd3281: Q <= 8'h02;
13'd3282: Q <= 8'h00;
13'd3283: Q <= 8'h00;
13'd3284: Q <= 8'h70;
13'd3285: Q <= 8'h50;
13'd3286: Q <= 8'h00;
13'd3287: Q <= 8'h00;
13'd3288: Q <= 8'h18;
13'd3289: Q <= 8'h50;
13'd3290: Q <= 8'h00;
13'd3291: Q <= 8'h00;
13'd3292: Q <= 8'hfd;
13'd3293: Q <= 8'h19;
13'd3294: Q <= 8'h11;
13'd3295: Q <= 8'h5d;
13'd3296: Q <= 8'h3f;
13'd3297: Q <= 8'h3b;
13'd3298: Q <= 8'h96;
13'd3299: Q <= 8'h4f;
13'd3300: Q <= 8'h40;
13'd3301: Q <= 8'hb5;
13'd3302: Q <= 8'ha4;
13'd3303: Q <= 8'h8a;
13'd3304: Q <= 8'h00;
13'd3305: Q <= 8'hcd;
13'd3306: Q <= 8'h50;
13'd3307: Q <= 8'h8c;
13'd3308: Q <= 8'h0e;
13'd3309: Q <= 8'hd5;
13'd3310: Q <= 8'h00;
13'd3311: Q <= 8'he0;
13'd3312: Q <= 8'h46;
13'd3313: Q <= 8'h5d;
13'd3314: Q <= 8'h14;
13'd3315: Q <= 8'h49;
13'd3316: Q <= 8'h0f;
13'd3317: Q <= 8'h5e;
13'd3318: Q <= 8'h07;
13'd3319: Q <= 8'h22;
13'd3320: Q <= 8'hc4;
13'd3321: Q <= 8'h53;
13'd3322: Q <= 8'hc2;
13'd3323: Q <= 8'he4;
13'd3324: Q <= 8'h44;
13'd3325: Q <= 8'he5;
13'd3326: Q <= 8'h64;
13'd3327: Q <= 8'hc4;
13'd3328: Q <= 8'hfe;
13'd3329: Q <= 8'hd0;
13'd3330: Q <= 8'h14;
13'd3331: Q <= 8'h51;
13'd3332: Q <= 8'h88;
13'd3333: Q <= 8'h51;
13'd3334: Q <= 8'h01;
13'd3335: Q <= 8'h76;
13'd3336: Q <= 8'hb0;
13'd3337: Q <= 8'h94;
13'd3338: Q <= 8'h01;
13'd3339: Q <= 8'h03;
13'd3340: Q <= 8'hc8;
13'd3341: Q <= 8'h85;
13'd3342: Q <= 8'h1c;
13'd3343: Q <= 8'h01;
13'd3344: Q <= 8'hbb;
13'd3345: Q <= 8'hc2;
13'd3346: Q <= 8'h4a;
13'd3347: Q <= 8'h24;
13'd3348: Q <= 8'h42;
13'd3349: Q <= 8'h01;
13'd3350: Q <= 8'h00;
13'd3351: Q <= 8'h30;
13'd3352: Q <= 8'hb3;
13'd3353: Q <= 8'h41;
13'd3354: Q <= 8'h0d;
13'd3355: Q <= 8'h10;
13'd3356: Q <= 8'h26;
13'd3357: Q <= 8'h38;
13'd3358: Q <= 8'h10;
13'd3359: Q <= 8'h01;
13'd3360: Q <= 8'h90;
13'd3361: Q <= 8'hb0;
13'd3362: Q <= 8'h0c;
13'd3363: Q <= 8'h85;
13'd3364: Q <= 8'h40;
13'd3365: Q <= 8'h40;
13'd3366: Q <= 8'h00;
13'd3367: Q <= 8'h00;
13'd3368: Q <= 8'h10;
13'd3369: Q <= 8'h30;
13'd3370: Q <= 8'h00;
13'd3371: Q <= 8'h4c;
13'd3372: Q <= 8'h15;
13'd3373: Q <= 8'h40;
13'd3374: Q <= 8'h00;
13'd3375: Q <= 8'h00;
13'd3376: Q <= 8'h10;
13'd3377: Q <= 8'hb1;
13'd3378: Q <= 8'h45;
13'd3379: Q <= 8'hfd;
13'd3380: Q <= 8'h00;
13'd3381: Q <= 8'h81;
13'd3382: Q <= 8'h00;
13'd3383: Q <= 8'h41;
13'd3384: Q <= 8'h00;
13'd3385: Q <= 8'hb3;
13'd3386: Q <= 8'h10;
13'd3387: Q <= 8'h2e;
13'd3388: Q <= 8'h41;
13'd3389: Q <= 8'h98;
13'd3390: Q <= 8'h00;
13'd3391: Q <= 8'h22;
13'd3392: Q <= 8'h14;
13'd3393: Q <= 8'h62;
13'd3394: Q <= 8'h00;
13'd3395: Q <= 8'h20;
13'd3396: Q <= 8'h00;
13'd3397: Q <= 8'h08;
13'd3398: Q <= 8'h94;
13'd3399: Q <= 8'hbf;
13'd3400: Q <= 8'haf;
13'd3401: Q <= 8'h8f;
13'd3402: Q <= 8'h00;
13'd3403: Q <= 8'h2c;
13'd3404: Q <= 8'h34;
13'd3405: Q <= 8'h09;
13'd3406: Q <= 8'h8c;
13'd3407: Q <= 8'h39;
13'd3408: Q <= 8'h60;
13'd3409: Q <= 8'h84;
13'd3410: Q <= 8'h24;
13'd3411: Q <= 8'h7c;
13'd3412: Q <= 8'h30;
13'd3413: Q <= 8'h1a;
13'd3414: Q <= 8'h0f;
13'd3415: Q <= 8'hb3;
13'd3416: Q <= 8'h29;
13'd3417: Q <= 8'had;
13'd3418: Q <= 8'h28;
13'd3419: Q <= 8'h89;
13'd3420: Q <= 8'h28;
13'd3421: Q <= 8'h06;
13'd3422: Q <= 8'h08;
13'd3423: Q <= 8'h3b;
13'd3424: Q <= 8'h30;
13'd3425: Q <= 8'h14;
13'd3426: Q <= 8'hd0;
13'd3427: Q <= 8'h30;
13'd3428: Q <= 8'hf4;
13'd3429: Q <= 8'h5e;
13'd3430: Q <= 8'hf1;
13'd3431: Q <= 8'hf5;
13'd3432: Q <= 8'hbb;
13'd3433: Q <= 8'h23;
13'd3434: Q <= 8'h80;
13'd3435: Q <= 8'h11;
13'd3436: Q <= 8'hc9;
13'd3437: Q <= 8'h3f;
13'd3438: Q <= 8'hb9;
13'd3439: Q <= 8'h04;
13'd3440: Q <= 8'h20;
13'd3441: Q <= 8'h71;
13'd3442: Q <= 8'h1c;
13'd3443: Q <= 8'hd8;
13'd3444: Q <= 8'h71;
13'd3445: Q <= 8'hbf;
13'd3446: Q <= 8'hf9;
13'd3447: Q <= 8'hda;
13'd3448: Q <= 8'hc8;
13'd3449: Q <= 8'h38;
13'd3450: Q <= 8'h3d;
13'd3451: Q <= 8'hbf;
13'd3452: Q <= 8'h34;
13'd3453: Q <= 8'h12;
13'd3454: Q <= 8'h28;
13'd3455: Q <= 8'ha8;
13'd3456: Q <= 8'hcf;
13'd3457: Q <= 8'h43;
13'd3458: Q <= 8'h1b;
13'd3459: Q <= 8'h04;
13'd3460: Q <= 8'h97;
13'd3461: Q <= 8'hfb;
13'd3462: Q <= 8'hff;
13'd3463: Q <= 8'h03;
13'd3464: Q <= 8'h66;
13'd3465: Q <= 8'hbf;
13'd3466: Q <= 8'h4c;
13'd3467: Q <= 8'h54;
13'd3468: Q <= 8'h87;
13'd3469: Q <= 8'hf5;
13'd3470: Q <= 8'h2a;
13'd3471: Q <= 8'h32;
13'd3472: Q <= 8'h0f;
13'd3473: Q <= 8'h0f;
13'd3474: Q <= 8'hf2;
13'd3475: Q <= 8'h24;
13'd3476: Q <= 8'he2;
13'd3477: Q <= 8'haf;
13'd3478: Q <= 8'h5e;
13'd3479: Q <= 8'h46;
13'd3480: Q <= 8'h44;
13'd3481: Q <= 8'hdd;
13'd3482: Q <= 8'h7d;
13'd3483: Q <= 8'h40;
13'd3484: Q <= 8'hc2;
13'd3485: Q <= 8'hfa;
13'd3486: Q <= 8'hd1;
13'd3487: Q <= 8'hc1;
13'd3488: Q <= 8'hd5;
13'd3489: Q <= 8'h01;
13'd3490: Q <= 8'h38;
13'd3491: Q <= 8'h03;
13'd3492: Q <= 8'h16;
13'd3493: Q <= 8'hef;
13'd3494: Q <= 8'h64;
13'd3495: Q <= 8'h20;
13'd3496: Q <= 8'hf5;
13'd3497: Q <= 8'h21;
13'd3498: Q <= 8'ha7;
13'd3499: Q <= 8'h7e;
13'd3500: Q <= 8'he1;
13'd3501: Q <= 8'hae;
13'd3502: Q <= 8'had;
13'd3503: Q <= 8'h55;
13'd3504: Q <= 8'h31;
13'd3505: Q <= 8'h2d;
13'd3506: Q <= 8'he4;
13'd3507: Q <= 8'h06;
13'd3508: Q <= 8'h7e;
13'd3509: Q <= 8'h44;
13'd3510: Q <= 8'h46;
13'd3511: Q <= 8'h47;
13'd3512: Q <= 8'h2d;
13'd3513: Q <= 8'h01;
13'd3514: Q <= 8'h54;
13'd3515: Q <= 8'h41;
13'd3516: Q <= 8'h7c;
13'd3517: Q <= 8'h04;
13'd3518: Q <= 8'h95;
13'd3519: Q <= 8'h7f;
13'd3520: Q <= 8'hfa;
13'd3521: Q <= 8'h10;
13'd3522: Q <= 8'h00;
13'd3523: Q <= 8'h04;
13'd3524: Q <= 8'h90;
13'd3525: Q <= 8'h50;
13'd3526: Q <= 8'h90;
13'd3527: Q <= 8'h88;
13'd3528: Q <= 8'hb8;
13'd3529: Q <= 8'h12;
13'd3530: Q <= 8'h02;
13'd3531: Q <= 8'h91;
13'd3532: Q <= 8'h1c;
13'd3533: Q <= 8'h04;
13'd3534: Q <= 8'h8c;
13'd3535: Q <= 8'hcd;
13'd3536: Q <= 8'hbf;
13'd3537: Q <= 8'h0a;
13'd3538: Q <= 8'h00;
13'd3539: Q <= 8'h00;
13'd3540: Q <= 8'ha6;
13'd3541: Q <= 8'h48;
13'd3542: Q <= 8'ha8;
13'd3543: Q <= 8'h88;
13'd3544: Q <= 8'hbf;
13'd3545: Q <= 8'h02;
13'd3546: Q <= 8'h48;
13'd3547: Q <= 8'h10;
13'd3548: Q <= 8'h8c;
13'd3549: Q <= 8'h50;
13'd3550: Q <= 8'h88;
13'd3551: Q <= 8'h8c;
13'd3552: Q <= 8'h6f;
13'd3553: Q <= 8'h6b;
13'd3554: Q <= 8'hb3;
13'd3555: Q <= 8'hb9;
13'd3556: Q <= 8'h2b;
13'd3557: Q <= 8'h2d;
13'd3558: Q <= 8'ha7;
13'd3559: Q <= 8'h04;
13'd3560: Q <= 8'h42;
13'd3561: Q <= 8'hee;
13'd3562: Q <= 8'h77;
13'd3563: Q <= 8'h24;
13'd3564: Q <= 8'h9a;
13'd3565: Q <= 8'h0c;
13'd3566: Q <= 8'h23;
13'd3567: Q <= 8'h20;
13'd3568: Q <= 8'h17;
13'd3569: Q <= 8'h0c;
13'd3570: Q <= 8'hda;
13'd3571: Q <= 8'h4c;
13'd3572: Q <= 8'hfb;
13'd3573: Q <= 8'h5c;
13'd3574: Q <= 8'h65;
13'd3575: Q <= 8'h62;
13'd3576: Q <= 8'h52;
13'd3577: Q <= 8'h16;
13'd3578: Q <= 8'h33;
13'd3579: Q <= 8'h35;
13'd3580: Q <= 8'h23;
13'd3581: Q <= 8'h37;
13'd3582: Q <= 8'h67;
13'd3583: Q <= 8'h55;
13'd3584: Q <= 8'h20;
13'd3585: Q <= 8'h00;
13'd3586: Q <= 8'h00;
13'd3587: Q <= 8'h11;
13'd3588: Q <= 8'h48;
13'd3589: Q <= 8'h10;
13'd3590: Q <= 8'had;
13'd3591: Q <= 8'h04;
13'd3592: Q <= 8'h3e;
13'd3593: Q <= 8'h00;
13'd3594: Q <= 8'h1d;
13'd3595: Q <= 8'h27;
13'd3596: Q <= 8'hbd;
13'd3597: Q <= 8'h15;
13'd3598: Q <= 8'hbd;
13'd3599: Q <= 8'h0f;
13'd3600: Q <= 8'ha0;
13'd3601: Q <= 8'h00;
13'd3602: Q <= 8'ha8;
13'd3603: Q <= 8'h01;
13'd3604: Q <= 8'h88;
13'd3605: Q <= 8'h90;
13'd3606: Q <= 8'h88;
13'd3607: Q <= 8'h4f;
13'd3608: Q <= 8'h84;
13'd3609: Q <= 8'hac;
13'd3610: Q <= 8'ha4;
13'd3611: Q <= 8'h20;
13'd3612: Q <= 8'hbb;
13'd3613: Q <= 8'h18;
13'd3614: Q <= 8'h18;
13'd3615: Q <= 8'h08;
13'd3616: Q <= 8'hcb;
13'd3617: Q <= 8'h93;
13'd3618: Q <= 8'h9f;
13'd3619: Q <= 8'heb;
13'd3620: Q <= 8'hff;
13'd3621: Q <= 8'hfe;
13'd3622: Q <= 8'hef;
13'd3623: Q <= 8'he7;
13'd3624: Q <= 8'h00;
13'd3625: Q <= 8'h50;
13'd3626: Q <= 8'hd1;
13'd3627: Q <= 8'h20;
13'd3628: Q <= 8'h12;
13'd3629: Q <= 8'hf8;
13'd3630: Q <= 8'h9e;
13'd3631: Q <= 8'ha0;
13'd3632: Q <= 8'h2e;
13'd3633: Q <= 8'h08;
13'd3634: Q <= 8'h6a;
13'd3635: Q <= 8'h40;
13'd3636: Q <= 8'h46;
13'd3637: Q <= 8'hf0;
13'd3638: Q <= 8'h4e;
13'd3639: Q <= 8'hc7;
13'd3640: Q <= 8'h54;
13'd3641: Q <= 8'h10;
13'd3642: Q <= 8'hc4;
13'd3643: Q <= 8'h52;
13'd3644: Q <= 8'he0;
13'd3645: Q <= 8'h54;
13'd3646: Q <= 8'hc4;
13'd3647: Q <= 8'h44;
13'd3648: Q <= 8'hbd;
13'd3649: Q <= 8'h16;
13'd3650: Q <= 8'hfb;
13'd3651: Q <= 8'h22;
13'd3652: Q <= 8'h17;
13'd3653: Q <= 8'h7b;
13'd3654: Q <= 8'h35;
13'd3655: Q <= 8'h0c;
13'd3656: Q <= 8'hf3;
13'd3657: Q <= 8'hb6;
13'd3658: Q <= 8'hff;
13'd3659: Q <= 8'h05;
13'd3660: Q <= 8'hfd;
13'd3661: Q <= 8'hf7;
13'd3662: Q <= 8'h57;
13'd3663: Q <= 8'h02;
13'd3664: Q <= 8'hc9;
13'd3665: Q <= 8'h84;
13'd3666: Q <= 8'hff;
13'd3667: Q <= 8'h46;
13'd3668: Q <= 8'h9e;
13'd3669: Q <= 8'hfc;
13'd3670: Q <= 8'hef;
13'd3671: Q <= 8'hd5;
13'd3672: Q <= 8'h8c;
13'd3673: Q <= 8'ha1;
13'd3674: Q <= 8'hbf;
13'd3675: Q <= 8'he4;
13'd3676: Q <= 8'hec;
13'd3677: Q <= 8'hb8;
13'd3678: Q <= 8'h84;
13'd3679: Q <= 8'h04;
13'd3680: Q <= 8'h35;
13'd3681: Q <= 8'h00;
13'd3682: Q <= 8'hd4;
13'd3683: Q <= 8'h18;
13'd3684: Q <= 8'hb5;
13'd3685: Q <= 8'h0d;
13'd3686: Q <= 8'h76;
13'd3687: Q <= 8'hdf;
13'd3688: Q <= 8'hdf;
13'd3689: Q <= 8'h17;
13'd3690: Q <= 8'h28;
13'd3691: Q <= 8'h28;
13'd3692: Q <= 8'h1d;
13'd3693: Q <= 8'h19;
13'd3694: Q <= 8'h3a;
13'd3695: Q <= 8'h2e;
13'd3696: Q <= 8'hbd;
13'd3697: Q <= 8'h0d;
13'd3698: Q <= 8'hbe;
13'd3699: Q <= 8'h0f;
13'd3700: Q <= 8'h5f;
13'd3701: Q <= 8'hdf;
13'd3702: Q <= 8'hfd;
13'd3703: Q <= 8'hff;
13'd3704: Q <= 8'hfd;
13'd3705: Q <= 8'h00;
13'd3706: Q <= 8'hee;
13'd3707: Q <= 8'h0a;
13'd3708: Q <= 8'h10;
13'd3709: Q <= 8'h09;
13'd3710: Q <= 8'h30;
13'd3711: Q <= 8'h0c;
13'd3712: Q <= 8'h3b;
13'd3713: Q <= 8'h39;
13'd3714: Q <= 8'h2f;
13'd3715: Q <= 8'h3d;
13'd3716: Q <= 8'hf9;
13'd3717: Q <= 8'hfc;
13'd3718: Q <= 8'h25;
13'd3719: Q <= 8'h23;
13'd3720: Q <= 8'he0;
13'd3721: Q <= 8'heb;
13'd3722: Q <= 8'hbd;
13'd3723: Q <= 8'h67;
13'd3724: Q <= 8'h80;
13'd3725: Q <= 8'h3e;
13'd3726: Q <= 8'h35;
13'd3727: Q <= 8'h5d;
13'd3728: Q <= 8'h01;
13'd3729: Q <= 8'ha9;
13'd3730: Q <= 8'h9f;
13'd3731: Q <= 8'haf;
13'd3732: Q <= 8'h38;
13'd3733: Q <= 8'h5f;
13'd3734: Q <= 8'h9e;
13'd3735: Q <= 8'h03;
13'd3736: Q <= 8'h30;
13'd3737: Q <= 8'h05;
13'd3738: Q <= 8'h27;
13'd3739: Q <= 8'h42;
13'd3740: Q <= 8'ha4;
13'd3741: Q <= 8'hb0;
13'd3742: Q <= 8'hc8;
13'd3743: Q <= 8'h25;
13'd3744: Q <= 8'h6f;
13'd3745: Q <= 8'h09;
13'd3746: Q <= 8'h5c;
13'd3747: Q <= 8'h56;
13'd3748: Q <= 8'h7f;
13'd3749: Q <= 8'h19;
13'd3750: Q <= 8'h7c;
13'd3751: Q <= 8'h1c;
13'd3752: Q <= 8'h4f;
13'd3753: Q <= 8'h16;
13'd3754: Q <= 8'h00;
13'd3755: Q <= 8'h6a;
13'd3756: Q <= 8'h4e;
13'd3757: Q <= 8'h2a;
13'd3758: Q <= 8'h0a;
13'd3759: Q <= 8'h2e;
13'd3760: Q <= 8'h57;
13'd3761: Q <= 8'h10;
13'd3762: Q <= 8'hb0;
13'd3763: Q <= 8'h6a;
13'd3764: Q <= 8'h5c;
13'd3765: Q <= 8'h0a;
13'd3766: Q <= 8'h16;
13'd3767: Q <= 8'h60;
13'd3768: Q <= 8'h44;
13'd3769: Q <= 8'h01;
13'd3770: Q <= 8'h00;
13'd3771: Q <= 8'h30;
13'd3772: Q <= 8'h40;
13'd3773: Q <= 8'h09;
13'd3774: Q <= 8'h64;
13'd3775: Q <= 8'h54;
13'd3776: Q <= 8'h6f;
13'd3777: Q <= 8'hdb;
13'd3778: Q <= 8'haf;
13'd3779: Q <= 8'he7;
13'd3780: Q <= 8'h43;
13'd3781: Q <= 8'h7b;
13'd3782: Q <= 8'hb7;
13'd3783: Q <= 8'h22;
13'd3784: Q <= 8'h60;
13'd3785: Q <= 8'h8d;
13'd3786: Q <= 8'hdc;
13'd3787: Q <= 8'hfc;
13'd3788: Q <= 8'h87;
13'd3789: Q <= 8'hc0;
13'd3790: Q <= 8'h13;
13'd3791: Q <= 8'h00;
13'd3792: Q <= 8'h6c;
13'd3793: Q <= 8'h56;
13'd3794: Q <= 8'hfe;
13'd3795: Q <= 8'h10;
13'd3796: Q <= 8'h2d;
13'd3797: Q <= 8'hcf;
13'd3798: Q <= 8'h72;
13'd3799: Q <= 8'h04;
13'd3800: Q <= 8'h54;
13'd3801: Q <= 8'h46;
13'd3802: Q <= 8'h72;
13'd3803: Q <= 8'h90;
13'd3804: Q <= 8'hf5;
13'd3805: Q <= 8'hdf;
13'd3806: Q <= 8'hf0;
13'd3807: Q <= 8'hc0;
13'd3808: Q <= 8'hef;
13'd3809: Q <= 8'hef;
13'd3810: Q <= 8'hff;
13'd3811: Q <= 8'hff;
13'd3812: Q <= 8'h30;
13'd3813: Q <= 8'h6b;
13'd3814: Q <= 8'h13;
13'd3815: Q <= 8'h4b;
13'd3816: Q <= 8'h43;
13'd3817: Q <= 8'h2e;
13'd3818: Q <= 8'h77;
13'd3819: Q <= 8'h32;
13'd3820: Q <= 8'h3b;
13'd3821: Q <= 8'ha6;
13'd3822: Q <= 8'h03;
13'd3823: Q <= 8'h06;
13'd3824: Q <= 8'h4b;
13'd3825: Q <= 8'hd7;
13'd3826: Q <= 8'h6f;
13'd3827: Q <= 8'h92;
13'd3828: Q <= 8'h17;
13'd3829: Q <= 8'h7f;
13'd3830: Q <= 8'h6b;
13'd3831: Q <= 8'h04;
13'd3832: Q <= 8'h23;
13'd3833: Q <= 8'h45;
13'd3834: Q <= 8'h67;
13'd3835: Q <= 8'h05;
13'd3836: Q <= 8'h57;
13'd3837: Q <= 8'hf7;
13'd3838: Q <= 8'h07;
13'd3839: Q <= 8'h40;
13'd3840: Q <= 8'h10;
13'd3841: Q <= 8'h10;
13'd3842: Q <= 8'h00;
13'd3843: Q <= 8'h11;
13'd3844: Q <= 8'h40;
13'd3845: Q <= 8'h24;
13'd3846: Q <= 8'h11;
13'd3847: Q <= 8'h31;
13'd3848: Q <= 8'h94;
13'd3849: Q <= 8'h90;
13'd3850: Q <= 8'h10;
13'd3851: Q <= 8'h00;
13'd3852: Q <= 8'h01;
13'd3853: Q <= 8'h80;
13'd3854: Q <= 8'h10;
13'd3855: Q <= 8'h00;
13'd3856: Q <= 8'h02;
13'd3857: Q <= 8'h01;
13'd3858: Q <= 8'h00;
13'd3859: Q <= 8'hb8;
13'd3860: Q <= 8'h90;
13'd3861: Q <= 8'h00;
13'd3862: Q <= 8'h08;
13'd3863: Q <= 8'hbb;
13'd3864: Q <= 8'h02;
13'd3865: Q <= 8'h48;
13'd3866: Q <= 8'h00;
13'd3867: Q <= 8'h83;
13'd3868: Q <= 8'h10;
13'd3869: Q <= 8'h00;
13'd3870: Q <= 8'h20;
13'd3871: Q <= 8'h00;
13'd3872: Q <= 8'hb0;
13'd3873: Q <= 8'h30;
13'd3874: Q <= 8'h00;
13'd3875: Q <= 8'h00;
13'd3876: Q <= 8'ha0;
13'd3877: Q <= 8'h10;
13'd3878: Q <= 8'h00;
13'd3879: Q <= 8'h20;
13'd3880: Q <= 8'ha0;
13'd3881: Q <= 8'h14;
13'd3882: Q <= 8'h00;
13'd3883: Q <= 8'h80;
13'd3884: Q <= 8'h80;
13'd3885: Q <= 8'h00;
13'd3886: Q <= 8'h00;
13'd3887: Q <= 8'h81;
13'd3888: Q <= 8'h73;
13'd3889: Q <= 8'h41;
13'd3890: Q <= 8'h40;
13'd3891: Q <= 8'h02;
13'd3892: Q <= 8'hb2;
13'd3893: Q <= 8'h02;
13'd3894: Q <= 8'ha0;
13'd3895: Q <= 8'h33;
13'd3896: Q <= 8'h77;
13'd3897: Q <= 8'h3b;
13'd3898: Q <= 8'h00;
13'd3899: Q <= 8'h13;
13'd3900: Q <= 8'h00;
13'd3901: Q <= 8'h01;
13'd3902: Q <= 8'h00;
13'd3903: Q <= 8'h53;
13'd3904: Q <= 8'hc0;
13'd3905: Q <= 8'h84;
13'd3906: Q <= 8'h00;
13'd3907: Q <= 8'h80;
13'd3908: Q <= 8'h04;
13'd3909: Q <= 8'h51;
13'd3910: Q <= 8'h00;
13'd3911: Q <= 8'h00;
13'd3912: Q <= 8'h84;
13'd3913: Q <= 8'h44;
13'd3914: Q <= 8'h00;
13'd3915: Q <= 8'h01;
13'd3916: Q <= 8'h05;
13'd3917: Q <= 8'h55;
13'd3918: Q <= 8'h04;
13'd3919: Q <= 8'h8c;
13'd3920: Q <= 8'h45;
13'd3921: Q <= 8'h41;
13'd3922: Q <= 8'h00;
13'd3923: Q <= 8'h00;
13'd3924: Q <= 8'h00;
13'd3925: Q <= 8'h00;
13'd3926: Q <= 8'h00;
13'd3927: Q <= 8'h00;
13'd3928: Q <= 8'h44;
13'd3929: Q <= 8'h45;
13'd3930: Q <= 8'h80;
13'd3931: Q <= 8'h00;
13'd3932: Q <= 8'hc0;
13'd3933: Q <= 8'h74;
13'd3934: Q <= 8'h08;
13'd3935: Q <= 8'h04;
13'd3936: Q <= 8'ha0;
13'd3937: Q <= 8'h09;
13'd3938: Q <= 8'h40;
13'd3939: Q <= 8'h09;
13'd3940: Q <= 8'h90;
13'd3941: Q <= 8'h19;
13'd3942: Q <= 8'h60;
13'd3943: Q <= 8'hcc;
13'd3944: Q <= 8'h84;
13'd3945: Q <= 8'h85;
13'd3946: Q <= 8'h91;
13'd3947: Q <= 8'h9d;
13'd3948: Q <= 8'h53;
13'd3949: Q <= 8'h05;
13'd3950: Q <= 8'h52;
13'd3951: Q <= 8'hdf;
13'd3952: Q <= 8'hbb;
13'd3953: Q <= 8'h08;
13'd3954: Q <= 8'h90;
13'd3955: Q <= 8'h1c;
13'd3956: Q <= 8'hf0;
13'd3957: Q <= 8'h01;
13'd3958: Q <= 8'hb0;
13'd3959: Q <= 8'h1a;
13'd3960: Q <= 8'hff;
13'd3961: Q <= 8'h18;
13'd3962: Q <= 8'h48;
13'd3963: Q <= 8'haf;
13'd3964: Q <= 8'h0c;
13'd3965: Q <= 8'h0a;
13'd3966: Q <= 8'h9c;
13'd3967: Q <= 8'h0f;
13'd3968: Q <= 8'hd1;
13'd3969: Q <= 8'h19;
13'd3970: Q <= 8'h6e;
13'd3971: Q <= 8'h0d;
13'd3972: Q <= 8'h10;
13'd3973: Q <= 8'h5d;
13'd3974: Q <= 8'h00;
13'd3975: Q <= 8'h0f;
13'd3976: Q <= 8'h71;
13'd3977: Q <= 8'h49;
13'd3978: Q <= 8'h5f;
13'd3979: Q <= 8'h1d;
13'd3980: Q <= 8'h10;
13'd3981: Q <= 8'h2d;
13'd3982: Q <= 8'h3a;
13'd3983: Q <= 8'h2f;
13'd3984: Q <= 8'hfe;
13'd3985: Q <= 8'h0d;
13'd3986: Q <= 8'hba;
13'd3987: Q <= 8'h4c;
13'd3988: Q <= 8'hbe;
13'd3989: Q <= 8'hae;
13'd3990: Q <= 8'hee;
13'd3991: Q <= 8'hac;
13'd3992: Q <= 8'hc5;
13'd3993: Q <= 8'h07;
13'd3994: Q <= 8'hac;
13'd3995: Q <= 8'h00;
13'd3996: Q <= 8'h10;
13'd3997: Q <= 8'h00;
13'd3998: Q <= 8'hc0;
13'd3999: Q <= 8'h0c;
13'd4000: Q <= 8'h59;
13'd4001: Q <= 8'h37;
13'd4002: Q <= 8'hc8;
13'd4003: Q <= 8'h16;
13'd4004: Q <= 8'h98;
13'd4005: Q <= 8'h34;
13'd4006: Q <= 8'h55;
13'd4007: Q <= 8'h77;
13'd4008: Q <= 8'hff;
13'd4009: Q <= 8'h5f;
13'd4010: Q <= 8'h10;
13'd4011: Q <= 8'h03;
13'd4012: Q <= 8'h15;
13'd4013: Q <= 8'h16;
13'd4014: Q <= 8'h20;
13'd4015: Q <= 8'h16;
13'd4016: Q <= 8'hfc;
13'd4017: Q <= 8'h07;
13'd4018: Q <= 8'h04;
13'd4019: Q <= 8'h37;
13'd4020: Q <= 8'h50;
13'd4021: Q <= 8'h1d;
13'd4022: Q <= 8'h46;
13'd4023: Q <= 8'h7f;
13'd4024: Q <= 8'ha6;
13'd4025: Q <= 8'h41;
13'd4026: Q <= 8'h26;
13'd4027: Q <= 8'h7b;
13'd4028: Q <= 8'h00;
13'd4029: Q <= 8'h2a;
13'd4030: Q <= 8'h24;
13'd4031: Q <= 8'h3e;
13'd4032: Q <= 8'ha3;
13'd4033: Q <= 8'ha8;
13'd4034: Q <= 8'h64;
13'd4035: Q <= 8'h25;
13'd4036: Q <= 8'hec;
13'd4037: Q <= 8'hec;
13'd4038: Q <= 8'he0;
13'd4039: Q <= 8'h02;
13'd4040: Q <= 8'h0f;
13'd4041: Q <= 8'hbe;
13'd4042: Q <= 8'hc0;
13'd4043: Q <= 8'ha1;
13'd4044: Q <= 8'h35;
13'd4045: Q <= 8'hc7;
13'd4046: Q <= 8'h00;
13'd4047: Q <= 8'h1a;
13'd4048: Q <= 8'h2b;
13'd4049: Q <= 8'h44;
13'd4050: Q <= 8'h46;
13'd4051: Q <= 8'h06;
13'd4052: Q <= 8'hc4;
13'd4053: Q <= 8'hfe;
13'd4054: Q <= 8'h95;
13'd4055: Q <= 8'h55;
13'd4056: Q <= 8'h27;
13'd4057: Q <= 8'h0b;
13'd4058: Q <= 8'h09;
13'd4059: Q <= 8'h26;
13'd4060: Q <= 8'hb5;
13'd4061: Q <= 8'h35;
13'd4062: Q <= 8'h3f;
13'd4063: Q <= 8'h3f;
13'd4064: Q <= 8'h4c;
13'd4065: Q <= 8'h29;
13'd4066: Q <= 8'h80;
13'd4067: Q <= 8'h00;
13'd4068: Q <= 8'hd4;
13'd4069: Q <= 8'h8e;
13'd4070: Q <= 8'hee;
13'd4071: Q <= 8'hc0;
13'd4072: Q <= 8'h1f;
13'd4073: Q <= 8'h0e;
13'd4074: Q <= 8'h04;
13'd4075: Q <= 8'h25;
13'd4076: Q <= 8'h4b;
13'd4077: Q <= 8'h02;
13'd4078: Q <= 8'hf6;
13'd4079: Q <= 8'h0e;
13'd4080: Q <= 8'h02;
13'd4081: Q <= 8'h00;
13'd4082: Q <= 8'hc0;
13'd4083: Q <= 8'h00;
13'd4084: Q <= 8'h5a;
13'd4085: Q <= 8'h00;
13'd4086: Q <= 8'h40;
13'd4087: Q <= 8'h22;
13'd4088: Q <= 8'h5c;
13'd4089: Q <= 8'h4e;
13'd4090: Q <= 8'h45;
13'd4091: Q <= 8'h3b;
13'd4092: Q <= 8'h24;
13'd4093: Q <= 8'h02;
13'd4094: Q <= 8'h40;
13'd4095: Q <= 8'h62;
13'd4096: Q <= 8'h03;
13'd4097: Q <= 8'h4e;
13'd4098: Q <= 8'hc3;
13'd4099: Q <= 8'h14;
13'd4100: Q <= 8'h0b;
13'd4101: Q <= 8'heb;
13'd4102: Q <= 8'h46;
13'd4103: Q <= 8'h40;
13'd4104: Q <= 8'h0a;
13'd4105: Q <= 8'h01;
13'd4106: Q <= 8'h9a;
13'd4107: Q <= 8'h99;
13'd4108: Q <= 8'h12;
13'd4109: Q <= 8'h92;
13'd4110: Q <= 8'h42;
13'd4111: Q <= 8'hea;
13'd4112: Q <= 8'h41;
13'd4113: Q <= 8'h43;
13'd4114: Q <= 8'h53;
13'd4115: Q <= 8'h6a;
13'd4116: Q <= 8'hc0;
13'd4117: Q <= 8'h82;
13'd4118: Q <= 8'h4a;
13'd4119: Q <= 8'h00;
13'd4120: Q <= 8'h01;
13'd4121: Q <= 8'h00;
13'd4122: Q <= 8'h46;
13'd4123: Q <= 8'h1b;
13'd4124: Q <= 8'h6f;
13'd4125: Q <= 8'hf5;
13'd4126: Q <= 8'h30;
13'd4127: Q <= 8'h40;
13'd4128: Q <= 8'h45;
13'd4129: Q <= 8'h75;
13'd4130: Q <= 8'hd1;
13'd4131: Q <= 8'h75;
13'd4132: Q <= 8'h63;
13'd4133: Q <= 8'he2;
13'd4134: Q <= 8'h29;
13'd4135: Q <= 8'h11;
13'd4136: Q <= 8'ha1;
13'd4137: Q <= 8'hea;
13'd4138: Q <= 8'he9;
13'd4139: Q <= 8'h62;
13'd4140: Q <= 8'hf3;
13'd4141: Q <= 8'hee;
13'd4142: Q <= 8'h0b;
13'd4143: Q <= 8'h00;
13'd4144: Q <= 8'h4e;
13'd4145: Q <= 8'hda;
13'd4146: Q <= 8'h66;
13'd4147: Q <= 8'hfd;
13'd4148: Q <= 8'hf7;
13'd4149: Q <= 8'hf6;
13'd4150: Q <= 8'h09;
13'd4151: Q <= 8'h1b;
13'd4152: Q <= 8'h4f;
13'd4153: Q <= 8'h77;
13'd4154: Q <= 8'h70;
13'd4155: Q <= 8'haa;
13'd4156: Q <= 8'h60;
13'd4157: Q <= 8'h68;
13'd4158: Q <= 8'h38;
13'd4159: Q <= 8'h40;
13'd4160: Q <= 8'h0c;
13'd4161: Q <= 8'h08;
13'd4162: Q <= 8'h00;
13'd4163: Q <= 8'h04;
13'd4164: Q <= 8'h9c;
13'd4165: Q <= 8'h06;
13'd4166: Q <= 8'h1d;
13'd4167: Q <= 8'hff;
13'd4168: Q <= 8'hcf;
13'd4169: Q <= 8'h68;
13'd4170: Q <= 8'h80;
13'd4171: Q <= 8'h08;
13'd4172: Q <= 8'h1f;
13'd4173: Q <= 8'h58;
13'd4174: Q <= 8'hce;
13'd4175: Q <= 8'h4f;
13'd4176: Q <= 8'h34;
13'd4177: Q <= 8'ha2;
13'd4178: Q <= 8'h01;
13'd4179: Q <= 8'h86;
13'd4180: Q <= 8'h0a;
13'd4181: Q <= 8'h28;
13'd4182: Q <= 8'h42;
13'd4183: Q <= 8'h7b;
13'd4184: Q <= 8'h1f;
13'd4185: Q <= 8'h1e;
13'd4186: Q <= 8'h2c;
13'd4187: Q <= 8'ha8;
13'd4188: Q <= 8'h3c;
13'd4189: Q <= 8'h08;
13'd4190: Q <= 8'h10;
13'd4191: Q <= 8'h2f;
13'd4192: Q <= 8'hdc;
13'd4193: Q <= 8'hd0;
13'd4194: Q <= 8'h42;
13'd4195: Q <= 8'h10;
13'd4196: Q <= 8'h70;
13'd4197: Q <= 8'h10;
13'd4198: Q <= 8'h18;
13'd4199: Q <= 8'h00;
13'd4200: Q <= 8'hdc;
13'd4201: Q <= 8'h11;
13'd4202: Q <= 8'h11;
13'd4203: Q <= 8'h00;
13'd4204: Q <= 8'h17;
13'd4205: Q <= 8'h50;
13'd4206: Q <= 8'h30;
13'd4207: Q <= 8'h12;
13'd4208: Q <= 8'h80;
13'd4209: Q <= 8'h0e;
13'd4210: Q <= 8'h10;
13'd4211: Q <= 8'h00;
13'd4212: Q <= 8'hfb;
13'd4213: Q <= 8'h18;
13'd4214: Q <= 8'h01;
13'd4215: Q <= 8'h40;
13'd4216: Q <= 8'h11;
13'd4217: Q <= 8'h0c;
13'd4218: Q <= 8'h20;
13'd4219: Q <= 8'h20;
13'd4220: Q <= 8'hdd;
13'd4221: Q <= 8'hd9;
13'd4222: Q <= 8'h30;
13'd4223: Q <= 8'h15;
13'd4224: Q <= 8'hb8;
13'd4225: Q <= 8'h08;
13'd4226: Q <= 8'h00;
13'd4227: Q <= 8'h00;
13'd4228: Q <= 8'he1;
13'd4229: Q <= 8'hcc;
13'd4230: Q <= 8'hc8;
13'd4231: Q <= 8'h0c;
13'd4232: Q <= 8'h45;
13'd4233: Q <= 8'h15;
13'd4234: Q <= 8'h19;
13'd4235: Q <= 8'h20;
13'd4236: Q <= 8'hc0;
13'd4237: Q <= 8'h50;
13'd4238: Q <= 8'hcd;
13'd4239: Q <= 8'hdd;
13'd4240: Q <= 8'hfa;
13'd4241: Q <= 8'h1c;
13'd4242: Q <= 8'h80;
13'd4243: Q <= 8'h09;
13'd4244: Q <= 8'hae;
13'd4245: Q <= 8'h88;
13'd4246: Q <= 8'h22;
13'd4247: Q <= 8'h89;
13'd4248: Q <= 8'h71;
13'd4249: Q <= 8'h10;
13'd4250: Q <= 8'h0a;
13'd4251: Q <= 8'h3a;
13'd4252: Q <= 8'h04;
13'd4253: Q <= 8'h01;
13'd4254: Q <= 8'h20;
13'd4255: Q <= 8'h0c;
13'd4256: Q <= 8'h07;
13'd4257: Q <= 8'h07;
13'd4258: Q <= 8'h8f;
13'd4259: Q <= 8'h0f;
13'd4260: Q <= 8'h12;
13'd4261: Q <= 8'hd3;
13'd4262: Q <= 8'h4b;
13'd4263: Q <= 8'h4f;
13'd4264: Q <= 8'h00;
13'd4265: Q <= 8'h04;
13'd4266: Q <= 8'h42;
13'd4267: Q <= 8'h26;
13'd4268: Q <= 8'h02;
13'd4269: Q <= 8'h01;
13'd4270: Q <= 8'ha2;
13'd4271: Q <= 8'hc2;
13'd4272: Q <= 8'h07;
13'd4273: Q <= 8'h04;
13'd4274: Q <= 8'hdf;
13'd4275: Q <= 8'h4d;
13'd4276: Q <= 8'h0d;
13'd4277: Q <= 8'hcb;
13'd4278: Q <= 8'h4b;
13'd4279: Q <= 8'h47;
13'd4280: Q <= 8'h61;
13'd4281: Q <= 8'h67;
13'd4282: Q <= 8'h2e;
13'd4283: Q <= 8'h5b;
13'd4284: Q <= 8'h10;
13'd4285: Q <= 8'h1d;
13'd4286: Q <= 8'h48;
13'd4287: Q <= 8'hd7;
13'd4288: Q <= 8'h47;
13'd4289: Q <= 8'h30;
13'd4290: Q <= 8'h27;
13'd4291: Q <= 8'h22;
13'd4292: Q <= 8'h03;
13'd4293: Q <= 8'h73;
13'd4294: Q <= 8'h07;
13'd4295: Q <= 8'h02;
13'd4296: Q <= 8'h48;
13'd4297: Q <= 8'h60;
13'd4298: Q <= 8'h06;
13'd4299: Q <= 8'h00;
13'd4300: Q <= 8'h04;
13'd4301: Q <= 8'hb2;
13'd4302: Q <= 8'h01;
13'd4303: Q <= 8'h00;
13'd4304: Q <= 8'h13;
13'd4305: Q <= 8'h6b;
13'd4306: Q <= 8'h6f;
13'd4307: Q <= 8'h55;
13'd4308: Q <= 8'h12;
13'd4309: Q <= 8'h30;
13'd4310: Q <= 8'h2f;
13'd4311: Q <= 8'h01;
13'd4312: Q <= 8'h57;
13'd4313: Q <= 8'h37;
13'd4314: Q <= 8'h7f;
13'd4315: Q <= 8'h72;
13'd4316: Q <= 8'h26;
13'd4317: Q <= 8'hf7;
13'd4318: Q <= 8'h42;
13'd4319: Q <= 8'h4c;
13'd4320: Q <= 8'h18;
13'd4321: Q <= 8'h33;
13'd4322: Q <= 8'h54;
13'd4323: Q <= 8'h25;
13'd4324: Q <= 8'ha0;
13'd4325: Q <= 8'h13;
13'd4326: Q <= 8'hac;
13'd4327: Q <= 8'h24;
13'd4328: Q <= 8'hdd;
13'd4329: Q <= 8'h4d;
13'd4330: Q <= 8'h89;
13'd4331: Q <= 8'h9d;
13'd4332: Q <= 8'h86;
13'd4333: Q <= 8'h15;
13'd4334: Q <= 8'hff;
13'd4335: Q <= 8'hcf;
13'd4336: Q <= 8'h8d;
13'd4337: Q <= 8'hbd;
13'd4338: Q <= 8'hcd;
13'd4339: Q <= 8'h87;
13'd4340: Q <= 8'hb0;
13'd4341: Q <= 8'h31;
13'd4342: Q <= 8'had;
13'd4343: Q <= 8'h19;
13'd4344: Q <= 8'h04;
13'd4345: Q <= 8'h05;
13'd4346: Q <= 8'had;
13'd4347: Q <= 8'h2f;
13'd4348: Q <= 8'h24;
13'd4349: Q <= 8'h00;
13'd4350: Q <= 8'hfd;
13'd4351: Q <= 8'h00;
13'd4352: Q <= 8'h0b;
13'd4353: Q <= 8'h6f;
13'd4354: Q <= 8'h3f;
13'd4355: Q <= 8'haf;
13'd4356: Q <= 8'h22;
13'd4357: Q <= 8'hb1;
13'd4358: Q <= 8'h06;
13'd4359: Q <= 8'h41;
13'd4360: Q <= 8'h21;
13'd4361: Q <= 8'h40;
13'd4362: Q <= 8'h32;
13'd4363: Q <= 8'h8a;
13'd4364: Q <= 8'h21;
13'd4365: Q <= 8'hf5;
13'd4366: Q <= 8'h04;
13'd4367: Q <= 8'h50;
13'd4368: Q <= 8'h63;
13'd4369: Q <= 8'h5a;
13'd4370: Q <= 8'h61;
13'd4371: Q <= 8'h6e;
13'd4372: Q <= 8'h14;
13'd4373: Q <= 8'hb7;
13'd4374: Q <= 8'h34;
13'd4375: Q <= 8'h47;
13'd4376: Q <= 8'h03;
13'd4377: Q <= 8'h58;
13'd4378: Q <= 8'hc1;
13'd4379: Q <= 8'h44;
13'd4380: Q <= 8'h71;
13'd4381: Q <= 8'hd5;
13'd4382: Q <= 8'h10;
13'd4383: Q <= 8'h42;
13'd4384: Q <= 8'hef;
13'd4385: Q <= 8'hfe;
13'd4386: Q <= 8'hef;
13'd4387: Q <= 8'hfb;
13'd4388: Q <= 8'h86;
13'd4389: Q <= 8'hfc;
13'd4390: Q <= 8'hcb;
13'd4391: Q <= 8'hb7;
13'd4392: Q <= 8'he2;
13'd4393: Q <= 8'h42;
13'd4394: Q <= 8'h2a;
13'd4395: Q <= 8'h12;
13'd4396: Q <= 8'h4f;
13'd4397: Q <= 8'ha5;
13'd4398: Q <= 8'ha3;
13'd4399: Q <= 8'hc0;
13'd4400: Q <= 8'h49;
13'd4401: Q <= 8'h50;
13'd4402: Q <= 8'h63;
13'd4403: Q <= 8'hd0;
13'd4404: Q <= 8'hc9;
13'd4405: Q <= 8'h00;
13'd4406: Q <= 8'h6c;
13'd4407: Q <= 8'h10;
13'd4408: Q <= 8'h44;
13'd4409: Q <= 8'hc0;
13'd4410: Q <= 8'h5d;
13'd4411: Q <= 8'hd9;
13'd4412: Q <= 8'h25;
13'd4413: Q <= 8'hc4;
13'd4414: Q <= 8'h44;
13'd4415: Q <= 8'h44;
13'd4416: Q <= 8'h9f;
13'd4417: Q <= 8'h27;
13'd4418: Q <= 8'h90;
13'd4419: Q <= 8'h20;
13'd4420: Q <= 8'h01;
13'd4421: Q <= 8'h00;
13'd4422: Q <= 8'h12;
13'd4423: Q <= 8'h61;
13'd4424: Q <= 8'h57;
13'd4425: Q <= 8'h00;
13'd4426: Q <= 8'hc0;
13'd4427: Q <= 8'h09;
13'd4428: Q <= 8'h41;
13'd4429: Q <= 8'h01;
13'd4430: Q <= 8'h02;
13'd4431: Q <= 8'h20;
13'd4432: Q <= 8'h04;
13'd4433: Q <= 8'h01;
13'd4434: Q <= 8'h83;
13'd4435: Q <= 8'h20;
13'd4436: Q <= 8'h2c;
13'd4437: Q <= 8'h00;
13'd4438: Q <= 8'h01;
13'd4439: Q <= 8'h4f;
13'd4440: Q <= 8'h0f;
13'd4441: Q <= 8'h28;
13'd4442: Q <= 8'had;
13'd4443: Q <= 8'h16;
13'd4444: Q <= 8'ha9;
13'd4445: Q <= 8'h05;
13'd4446: Q <= 8'h17;
13'd4447: Q <= 8'h3f;
        default: Q <= 0;
      endcase
    end
  end

endmodule

