module M_1
(
  output reg [40-1:0] Q,
  input wire [8-1:0] A,
  input wire cen,
  input wire clk,
  input wire reset

);

  always@(posedge clk) begin
    if(reset) begin
      Q <= 0;
    end
    else if(cen) begin
      case(A)
        //32'd0: Q <= 1;
        8'd0: Q <= 40'h1851030000;
8'd1: Q <= 40'h0471040000;
8'd2: Q <= 40'h0001830000;
8'd3: Q <= 40'h2c50c37230;
8'd4: Q <= 40'h0831046f21;
8'd5: Q <= 40'h3470c56656;
8'd6: Q <= 40'h18610474b0;
8'd7: Q <= 40'h18610269c0;
8'd8: Q <= 40'h0430c15fd7;
8'd9: Q <= 40'h0c11c361fa;
8'd10: Q <= 40'h00c20462c0;
8'd11: Q <= 40'h30210160f4;
8'd12: Q <= 40'h1060855d9f;
8'd13: Q <= 40'h2050c25ab2;
8'd14: Q <= 40'h3cd0c25618;
8'd15: Q <= 40'h1c91415e30;
8'd16: Q <= 40'h2401435838;
8'd17: Q <= 40'h00b0c453a7;
8'd18: Q <= 40'h3070c45472;
8'd19: Q <= 40'h1850835a74;
8'd20: Q <= 40'h0910c2555e;
8'd21: Q <= 40'h18310456ee;
8'd22: Q <= 40'h0040c3570b;
8'd23: Q <= 40'h24208650c6;
8'd24: Q <= 40'h3c60c251da;
8'd25: Q <= 40'h00e103517c;
8'd26: Q <= 40'h3460854eba;
8'd27: Q <= 40'h1000834c0f;
8'd28: Q <= 40'h1081034a1e;
8'd29: Q <= 40'h3c008264f6;
8'd30: Q <= 40'h2c308252d6;
8'd31: Q <= 40'h1c408354ea;
8'd32: Q <= 40'h30a0c24c6f;
8'd33: Q <= 40'h0800834efa;
8'd34: Q <= 40'h3520825594;
8'd35: Q <= 40'h2d10414c0c;
8'd36: Q <= 40'h1c00c74aaa;
8'd37: Q <= 40'h0c70844a60;
8'd38: Q <= 40'h3800824b27;
8'd39: Q <= 40'h2850c34b86;
8'd40: Q <= 40'h0810825164;
8'd41: Q <= 40'h28a0414c94;
8'd42: Q <= 40'h3d10824cb0;
8'd43: Q <= 40'h185085487a;
8'd44: Q <= 40'h3820c249c4;
8'd45: Q <= 40'h303043465f;
8'd46: Q <= 40'h0c00824808;
8'd47: Q <= 40'h1071424716;
8'd48: Q <= 40'h44c08246f0;
8'd49: Q <= 40'h04e10347c6;
8'd50: Q <= 40'h28a04248b6;
8'd51: Q <= 40'h38104346fa;
8'd52: Q <= 40'h35204246eb;
8'd53: Q <= 40'h14008245b6;
8'd54: Q <= 40'h14a0824a3a;
8'd55: Q <= 40'h38d0c34756;
8'd56: Q <= 40'h250081471c;
8'd57: Q <= 40'h2050824a54;
8'd58: Q <= 40'h08210645f0;
8'd59: Q <= 40'h04d1014681;
8'd60: Q <= 40'h4030844746;
8'd61: Q <= 40'h30e10349e8;
8'd62: Q <= 40'h2c8042439a;
8'd63: Q <= 40'h2120424508;
8'd64: Q <= 40'h0c7081446c;
8'd65: Q <= 40'h0d2082422c;
8'd66: Q <= 40'h401083431d;
8'd67: Q <= 40'h28704545aa;
8'd68: Q <= 40'h0010c33e20;
8'd69: Q <= 40'h28f0414144;
8'd70: Q <= 40'h3cb0c44578;
8'd71: Q <= 40'h1d5081409c;
8'd72: Q <= 40'h30108542a4;
8'd73: Q <= 40'h14608540b8;
8'd74: Q <= 40'h3c00834153;
8'd75: Q <= 40'h2ca041482a;
8'd76: Q <= 40'h04c0825174;
8'd77: Q <= 40'h2520414226;
8'd78: Q <= 40'h2c604140c8;
8'd79: Q <= 40'h291041400e;
8'd80: Q <= 40'h28e0c33f94;
8'd81: Q <= 40'h2000443fa4;
8'd82: Q <= 40'h28804142fe;
8'd83: Q <= 40'h1030814217;
8'd84: Q <= 40'h1490823eea;
8'd85: Q <= 40'h3510c24044;
8'd86: Q <= 40'h4060414144;
8'd87: Q <= 40'h251041406a;
8'd88: Q <= 40'h1920423f26;
8'd89: Q <= 40'h4410853fe2;
8'd90: Q <= 40'h0000c5400e;
8'd91: Q <= 40'h311041407e;
8'd92: Q <= 40'h1841034068;
8'd93: Q <= 40'h2ca042401f;
8'd94: Q <= 40'h3150814012;
8'd95: Q <= 40'h2c5106421c;
8'd96: Q <= 40'h0910c24262;
8'd97: Q <= 40'h2900414078;
8'd98: Q <= 40'h0010c73d20;
8'd99: Q <= 40'h0410823e86;
8'd100: Q <= 40'h1060813d7e;
8'd101: Q <= 40'h3c40c63e66;
8'd102: Q <= 40'h2850423d05;
8'd103: Q <= 40'h2110c13e9e;
8'd104: Q <= 40'h300082469c;
8'd105: Q <= 40'h2c70823d90;
8'd106: Q <= 40'h3d10c23e9c;
8'd107: Q <= 40'h0010833f5e;
8'd108: Q <= 40'h2900813e2a;
8'd109: Q <= 40'h38d0813e56;
8'd110: Q <= 40'h4410823e3e;
8'd111: Q <= 40'h2450414089;
8'd112: Q <= 40'h08b0833fa8;
8'd113: Q <= 40'h28f0813c38;
8'd114: Q <= 40'h0870813cd4;
8'd115: Q <= 40'h2890413b5a;
8'd116: Q <= 40'h1950813cca;
8'd117: Q <= 40'h3510823e6a;
8'd118: Q <= 40'h2d10413d5e;
8'd119: Q <= 40'h2950413e8e;
8'd120: Q <= 40'h0001023d99;
8'd121: Q <= 40'h3c40c23e0e;
8'd122: Q <= 40'h1431043ea4;
8'd123: Q <= 40'h0510c23f0a;
8'd124: Q <= 40'h30b0413faa;
8'd125: Q <= 40'h24b0413caa;
8'd126: Q <= 40'h30c0c23bea;
8'd127: Q <= 40'h3910823cf2;
8'd128: Q <= 40'h2d10413b84;
8'd129: Q <= 40'h0401434012;
8'd130: Q <= 40'h4100823ed1;
8'd131: Q <= 40'h2c50423e66;
8'd132: Q <= 40'h4800824556;
8'd133: Q <= 40'h38708139fe;
8'd134: Q <= 40'h2500413b0e;
8'd135: Q <= 40'h1120823c6a;
8'd136: Q <= 40'h2d20413ca4;
8'd137: Q <= 40'h2cf0413cca;
8'd138: Q <= 40'h34b0c23d4e;
8'd139: Q <= 40'h0000413cca;
8'd140: Q <= 40'h0000413d93;
8'd141: Q <= 40'h000041408c;
        default: Q <= 0;
      endcase
    end
  end

endmodule

