`define IN_NBYTE 1
`define PX_BLANKING 180
`define II_BIT_WIDTH 32
`define WIN_H 24
`define CLK_PERIOD 34
`define SIM_FRAMES 1
`define WIN_W 25
`define LOG_MAX_FDCNT 5
`define LOG_WIN_SIZE 10
`define LOG_NST 5
`define LOG_WIN_W 6
`define LOG_WIN_H 6
`define OUT_NBYTE 1
`define INIT_SCALE 0
`define SQII_BIT_WIDTH 32
`define WIN_SIZE 600
`define MAX_FDCNT 26
`define MAX_FRAME_W 320
`define NNVAR_BIT_WIDTH 32
`define HITVAL_ALL_PASS 100
`define LOG_MIN_LB_SIZE 13
`define SIZE 256
`define LOG_SIZE 8
`define SIM_TIME_LIMIT -1
`define HITVAL_FILLING 101
`define IM_SIZE 4096
`define LOG_IM_SIZE 12
`define LOG_FRAME_W 9
